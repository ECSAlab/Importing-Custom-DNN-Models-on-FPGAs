------------------------------------------HEADER START"------------------------------------------
--THIS FILE WAS GENERATED USING HIGH LANGUAGE DESCRIPTION TOOL DESIGNED BY: MUHAMMAD HAMDAN
--TOOL VERSION: 0.1
--GENERATION DATE/TIME:Tue Feb 09 00:01:34 CET 2021
------------------------------------------HEADER END"--------------------------------------------



------------------------------DESCRIPTION AND LIBRARY DECLARATION-START---------------------------
-- Engineer:       Muhammad Hamdan
-- Design Name:    HDL GENERATION - CONV LAYER 
-- Module Name:    FC - Behavioral 
-- Project Name:   CNN accelerator
-- Number of Total Operaiton: 40
-- Number of Clock Cycles: 48
-- Number of GOPS = 0.0
-------------------------------------------------Total Number of Operations for the Entire Model:10
-- Target Devices: Zynq-XC7Z020
-- Description: 
-- Dependencies: 
-- Revision:0.010 


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_arith.all;

entity FC_LAYER_7 is

GENERIC
 	( 
	constant PRECISION      : positive := 5; 	
	constant WHOLE          : positive := 2; 	
	constant DECIMAL        : positive := 3; 	
	constant DOUT_WIDTH     : positive := 5; 	
	constant BIAS_SIZE      : positive := 5;
	constant MULT_SIZE      : positive := 10;
	constant BASE_DIN_WIDTH : positive := 5;
	constant DIN_WIDTH      : positive := 5;
	constant IMAGE_WIDTH    : positive := 1;
	constant IMAGE_SIZE     : positive := 1024;	
	constant F_SIZE         : positive := 1;
	constant PF_X2_SIZE     : positive := 25;
	constant WEIGHT_SIZE    : positive := 5;
	constant BIASES_SIZE	: positive := 2;
	constant PADDING        : positive := 1;
	constant STRIDE         : positive := 1;
	constant FEATURE_MAPS   : positive := 10;
	constant VALID_CYCLES   : positive := 25;
	constant VALID_LOCAL_PIX: positive := 5;
	constant ADD_TREE_DEPTH : positive := 1;
	constant INPUT_DEPTH    : positive := 7;
	constant INNER_PXL_SUM  : positive := 1;
	constant SUM_PEXILS     : positive := 30;
	constant MULT_SUM_D_1   : positive := 60;
	constant MULT_SUM_SIZE_1: positive := 6;
	constant MULT_SUM_D_2   : positive := 30;
	constant MULT_SUM_SIZE_2: positive := 6;
	constant MULT_SUM_D_3   : positive := 15;
	constant MULT_SUM_SIZE_3: positive := 6;
	constant MULT_SUM_D_4   : positive := 8;
	constant MULT_SUM_SIZE_4: positive := 6;
	constant MULT_SUM_D_5   : positive := 4;
	constant MULT_SUM_SIZE_5: positive := 6;
	constant MULT_SUM_D_6   : positive := 2;
	constant MULT_SUM_SIZE_6: positive := 6;
	constant MULT_SUM_D_7   : positive := 1;
	constant MULT_SUM_SIZE_7: positive := 6;
	constant LOCAL_OUTPUT   : positive := 5	
		); 

port(
	DIN_1_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_2_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_3_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_4_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_5_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_6_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_7_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_8_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_9_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_10_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_11_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_12_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_13_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_14_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_15_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_16_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_17_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_18_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_19_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_20_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_21_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_22_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_23_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_24_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_25_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_26_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_27_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_28_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_29_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_30_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_31_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_32_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_33_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_34_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_35_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_36_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_37_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_38_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_39_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_40_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_41_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_42_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_43_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_44_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_45_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_46_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_47_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_48_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_49_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_50_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_51_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_52_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_53_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_54_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_55_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_56_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_57_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_58_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_59_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_60_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_61_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_62_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_63_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_64_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_65_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_66_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_67_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_68_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_69_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_70_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_71_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_72_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_73_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_74_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_75_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_76_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_77_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_78_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_79_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_80_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_81_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_82_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_83_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_84_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_85_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_86_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_87_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_88_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_89_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_90_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_91_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_92_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_93_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_94_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_95_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_96_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_97_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_98_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_99_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_100_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_101_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_102_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_103_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_104_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_105_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_106_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_107_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_108_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_109_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_110_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_111_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_112_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_113_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_114_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_115_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_116_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_117_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_118_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_119_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	DIN_120_7         :IN std_logic_vector(DIN_WIDTH-1 downto 0);
	CLK,RST         :IN std_logic;
   	DIS_STREAM      :OUT std_logic; 				-- S_AXIS_TVALID  : Data in is valid
   	EN_STREAM       :IN std_logic; 					-- S_AXIS_TREADY  : Ready to accept data in 
	EN_STREAM_OUT_7 :OUT std_logic; 			-- M_AXIS_TREADY  : Connected slave device is ready to accept data out/ Internal Enable
	VALID_OUT_7     :OUT std_logic;                         -- M_AXIS_TVALID  : Data out is valid
	EN_LOC_STREAM_7 :IN std_logic;
	DOUT_1_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_2_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_3_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_4_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_5_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_6_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_7_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_8_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_9_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	DOUT_10_7        :OUT std_logic_vector(DOUT_WIDTH-1 downto 0);
	INTERNAL_RST    :OUT std_logic
	);	

end FC_LAYER_7;

------------------------------ ARCHITECTURE DECLARATION - START---------------------------------------------

architecture Behavioral of FC_LAYER_7 is

------------------------------ INTERNAL FIXED CONSTANT & SIGNALS DECLARATION - START---------------------------------------------
type       FILTER_TYPE             is array (0 to PF_X2_SIZE-1) of signed(WEIGHT_SIZE- 1 downto 0);
signal     VALID_NXTLYR_PIX        :integer range 0 to VALID_CYCLES;
signal     PIXEL_COUNT             :integer range 0 to VALID_CYCLES;
signal     OUT_PIXEL_COUNT         :integer range 0 to VALID_CYCLES;
signal     EN_NXT_LYR_7            :std_logic;
signal     FRST_TIM_EN_7           :std_logic;
signal     Enable_MULT             :std_logic;
signal     Enable_ADDER            :std_logic;
signal     Enable_ReLU             :std_logic;
signal     Enable_BIAS             :std_logic;
signal     COUNT_PIX               :integer range 0 to PF_X2_SIZE;
signal     SIG_STRIDE              :integer range 0 to IMAGE_SIZE;
signal     PADDING_count           :integer range 0 to IMAGE_SIZE; -- TEMPORARY
signal     ROW_COUNT               :integer range 0 to IMAGE_SIZE; -- TEMPORARY


------------------------------ INTERNAL DYNAMIC SIGNALS DECLARATION ARRAY TYPE- START---------------------------------------------


type   MULT_X		is array (0 to FEATURE_MAPS-1) of signed(MULT_SIZE-1 downto 0);
signal MULT_1:MULT_X;
signal MULT_2:MULT_X;
signal MULT_3:MULT_X;
signal MULT_4:MULT_X;
signal MULT_5:MULT_X;
signal MULT_6:MULT_X;
signal MULT_7:MULT_X;
signal MULT_8:MULT_X;
signal MULT_9:MULT_X;
signal MULT_10:MULT_X;
signal MULT_11:MULT_X;
signal MULT_12:MULT_X;
signal MULT_13:MULT_X;
signal MULT_14:MULT_X;
signal MULT_15:MULT_X;
signal MULT_16:MULT_X;
signal MULT_17:MULT_X;
signal MULT_18:MULT_X;
signal MULT_19:MULT_X;
signal MULT_20:MULT_X;
signal MULT_21:MULT_X;
signal MULT_22:MULT_X;
signal MULT_23:MULT_X;
signal MULT_24:MULT_X;
signal MULT_25:MULT_X;
signal MULT_26:MULT_X;
signal MULT_27:MULT_X;
signal MULT_28:MULT_X;
signal MULT_29:MULT_X;
signal MULT_30:MULT_X;
signal MULT_31:MULT_X;
signal MULT_32:MULT_X;
signal MULT_33:MULT_X;
signal MULT_34:MULT_X;
signal MULT_35:MULT_X;
signal MULT_36:MULT_X;
signal MULT_37:MULT_X;
signal MULT_38:MULT_X;
signal MULT_39:MULT_X;
signal MULT_40:MULT_X;
signal MULT_41:MULT_X;
signal MULT_42:MULT_X;
signal MULT_43:MULT_X;
signal MULT_44:MULT_X;
signal MULT_45:MULT_X;
signal MULT_46:MULT_X;
signal MULT_47:MULT_X;
signal MULT_48:MULT_X;
signal MULT_49:MULT_X;
signal MULT_50:MULT_X;
signal MULT_51:MULT_X;
signal MULT_52:MULT_X;
signal MULT_53:MULT_X;
signal MULT_54:MULT_X;
signal MULT_55:MULT_X;
signal MULT_56:MULT_X;
signal MULT_57:MULT_X;
signal MULT_58:MULT_X;
signal MULT_59:MULT_X;
signal MULT_60:MULT_X;
signal MULT_61:MULT_X;
signal MULT_62:MULT_X;
signal MULT_63:MULT_X;
signal MULT_64:MULT_X;
signal MULT_65:MULT_X;
signal MULT_66:MULT_X;
signal MULT_67:MULT_X;
signal MULT_68:MULT_X;
signal MULT_69:MULT_X;
signal MULT_70:MULT_X;
signal MULT_71:MULT_X;
signal MULT_72:MULT_X;
signal MULT_73:MULT_X;
signal MULT_74:MULT_X;
signal MULT_75:MULT_X;
signal MULT_76:MULT_X;
signal MULT_77:MULT_X;
signal MULT_78:MULT_X;
signal MULT_79:MULT_X;
signal MULT_80:MULT_X;
signal MULT_81:MULT_X;
signal MULT_82:MULT_X;
signal MULT_83:MULT_X;
signal MULT_84:MULT_X;
signal MULT_85:MULT_X;
signal MULT_86:MULT_X;
signal MULT_87:MULT_X;
signal MULT_88:MULT_X;
signal MULT_89:MULT_X;
signal MULT_90:MULT_X;
signal MULT_91:MULT_X;
signal MULT_92:MULT_X;
signal MULT_93:MULT_X;
signal MULT_94:MULT_X;
signal MULT_95:MULT_X;
signal MULT_96:MULT_X;
signal MULT_97:MULT_X;
signal MULT_98:MULT_X;
signal MULT_99:MULT_X;
signal MULT_100:MULT_X;
signal MULT_101:MULT_X;
signal MULT_102:MULT_X;
signal MULT_103:MULT_X;
signal MULT_104:MULT_X;
signal MULT_105:MULT_X;
signal MULT_106:MULT_X;
signal MULT_107:MULT_X;
signal MULT_108:MULT_X;
signal MULT_109:MULT_X;
signal MULT_110:MULT_X;
signal MULT_111:MULT_X;
signal MULT_112:MULT_X;
signal MULT_113:MULT_X;
signal MULT_114:MULT_X;
signal MULT_115:MULT_X;
signal MULT_116:MULT_X;
signal MULT_117:MULT_X;
signal MULT_118:MULT_X;
signal MULT_119:MULT_X;
signal MULT_120:MULT_X;
signal DOUT_BUF_1_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_1		: signed(PRECISION-1 downto 0);
signal ReLU_1		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_2_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_2		: signed(PRECISION-1 downto 0);
signal ReLU_2		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_3_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_3		: signed(PRECISION-1 downto 0);
signal ReLU_3		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_4_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_4		: signed(PRECISION-1 downto 0);
signal ReLU_4		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_5_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_5		: signed(PRECISION-1 downto 0);
signal ReLU_5		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_6_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_6		: signed(PRECISION-1 downto 0);
signal ReLU_6		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_7_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_7		: signed(PRECISION-1 downto 0);
signal ReLU_7		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_8_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_8		: signed(PRECISION-1 downto 0);
signal ReLU_8		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_9_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_9		: signed(PRECISION-1 downto 0);
signal ReLU_9		: signed(PRECISION-1 downto 0);
signal DOUT_BUF_10_7	: std_logic_vector(LOCAL_OUTPUT-1 downto 0);
signal BIAS_10		: signed(PRECISION-1 downto 0);
signal ReLU_10		: signed(PRECISION-1 downto 0);


------------------------------------------------------ MULT SUMMATION DECLARATION-----------------------------------------------------------
signal SUM_PIXELS_1: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_2: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_3: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_4: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_5: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_6: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_7: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_8: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_9: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_10: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_11: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_12: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_13: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_14: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_15: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_16: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_17: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_18: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_19: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_20: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_21: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_22: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_23: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_24: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_25: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_26: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_27: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_28: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_29: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_30: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_31: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_32: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_33: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_34: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_35: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_36: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_37: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_38: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_39: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_40: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_41: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_42: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_43: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_44: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_45: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_46: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_47: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_48: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_49: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_50: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_51: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_52: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_53: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_54: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_55: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_56: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_57: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_58: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_59: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_60: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_61: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_62: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_63: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_64: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_65: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_66: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_67: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_68: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_69: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_70: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_71: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_72: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_73: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_74: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_75: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_76: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_77: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_78: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_79: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_80: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_81: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_82: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_83: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_84: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_85: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_86: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_87: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_88: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_89: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_90: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_91: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_92: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_93: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_94: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_95: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_96: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_97: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_98: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_99: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_100: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_101: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_102: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_103: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_104: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_105: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_106: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_107: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_108: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_109: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_110: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_111: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_112: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_113: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_114: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_115: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_116: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_117: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_118: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_119: signed(PRECISION-1 downto 0);
signal SUM_PIXELS_120: signed(PRECISION-1 downto 0);
type    MULT_X_SUM_1	is array (0 to FEATURE_MAPS-1) of signed(PRECISION-1 downto 0);
signal  EN_SUM_MULT_1	: std_logic;
signal  MULTS_1_1:MULT_X_SUM_1;
signal  MULTS_1_2:MULT_X_SUM_1;
signal  MULTS_1_3:MULT_X_SUM_1;
signal  MULTS_1_4:MULT_X_SUM_1;
signal  MULTS_1_5:MULT_X_SUM_1;
signal  MULTS_1_6:MULT_X_SUM_1;
signal  MULTS_1_7:MULT_X_SUM_1;
signal  MULTS_1_8:MULT_X_SUM_1;
signal  MULTS_1_9:MULT_X_SUM_1;
signal  MULTS_1_10:MULT_X_SUM_1;
signal  MULTS_1_11:MULT_X_SUM_1;
signal  MULTS_1_12:MULT_X_SUM_1;
signal  MULTS_1_13:MULT_X_SUM_1;
signal  MULTS_1_14:MULT_X_SUM_1;
signal  MULTS_1_15:MULT_X_SUM_1;
signal  MULTS_1_16:MULT_X_SUM_1;
signal  MULTS_1_17:MULT_X_SUM_1;
signal  MULTS_1_18:MULT_X_SUM_1;
signal  MULTS_1_19:MULT_X_SUM_1;
signal  MULTS_1_20:MULT_X_SUM_1;
signal  MULTS_1_21:MULT_X_SUM_1;
signal  MULTS_1_22:MULT_X_SUM_1;
signal  MULTS_1_23:MULT_X_SUM_1;
signal  MULTS_1_24:MULT_X_SUM_1;
signal  MULTS_1_25:MULT_X_SUM_1;
signal  MULTS_1_26:MULT_X_SUM_1;
signal  MULTS_1_27:MULT_X_SUM_1;
signal  MULTS_1_28:MULT_X_SUM_1;
signal  MULTS_1_29:MULT_X_SUM_1;
signal  MULTS_1_30:MULT_X_SUM_1;
signal  MULTS_1_31:MULT_X_SUM_1;
signal  MULTS_1_32:MULT_X_SUM_1;
signal  MULTS_1_33:MULT_X_SUM_1;
signal  MULTS_1_34:MULT_X_SUM_1;
signal  MULTS_1_35:MULT_X_SUM_1;
signal  MULTS_1_36:MULT_X_SUM_1;
signal  MULTS_1_37:MULT_X_SUM_1;
signal  MULTS_1_38:MULT_X_SUM_1;
signal  MULTS_1_39:MULT_X_SUM_1;
signal  MULTS_1_40:MULT_X_SUM_1;
signal  MULTS_1_41:MULT_X_SUM_1;
signal  MULTS_1_42:MULT_X_SUM_1;
signal  MULTS_1_43:MULT_X_SUM_1;
signal  MULTS_1_44:MULT_X_SUM_1;
signal  MULTS_1_45:MULT_X_SUM_1;
signal  MULTS_1_46:MULT_X_SUM_1;
signal  MULTS_1_47:MULT_X_SUM_1;
signal  MULTS_1_48:MULT_X_SUM_1;
signal  MULTS_1_49:MULT_X_SUM_1;
signal  MULTS_1_50:MULT_X_SUM_1;
signal  MULTS_1_51:MULT_X_SUM_1;
signal  MULTS_1_52:MULT_X_SUM_1;
signal  MULTS_1_53:MULT_X_SUM_1;
signal  MULTS_1_54:MULT_X_SUM_1;
signal  MULTS_1_55:MULT_X_SUM_1;
signal  MULTS_1_56:MULT_X_SUM_1;
signal  MULTS_1_57:MULT_X_SUM_1;
signal  MULTS_1_58:MULT_X_SUM_1;
signal  MULTS_1_59:MULT_X_SUM_1;
signal  MULTS_1_60:MULT_X_SUM_1;
signal  MULTS_1_61:MULT_X_SUM_1;
signal  MULTS_1_62:MULT_X_SUM_1;
signal  MULTS_1_63:MULT_X_SUM_1;
signal  MULTS_1_64:MULT_X_SUM_1;
signal  MULTS_1_65:MULT_X_SUM_1;
signal  MULTS_1_66:MULT_X_SUM_1;
signal  MULTS_1_67:MULT_X_SUM_1;
signal  MULTS_1_68:MULT_X_SUM_1;
signal  MULTS_1_69:MULT_X_SUM_1;
signal  MULTS_1_70:MULT_X_SUM_1;
signal  MULTS_1_71:MULT_X_SUM_1;
signal  MULTS_1_72:MULT_X_SUM_1;
signal  MULTS_1_73:MULT_X_SUM_1;
signal  MULTS_1_74:MULT_X_SUM_1;
signal  MULTS_1_75:MULT_X_SUM_1;
signal  MULTS_1_76:MULT_X_SUM_1;
signal  MULTS_1_77:MULT_X_SUM_1;
signal  MULTS_1_78:MULT_X_SUM_1;
signal  MULTS_1_79:MULT_X_SUM_1;
signal  MULTS_1_80:MULT_X_SUM_1;
signal  MULTS_1_81:MULT_X_SUM_1;
signal  MULTS_1_82:MULT_X_SUM_1;
signal  MULTS_1_83:MULT_X_SUM_1;
signal  MULTS_1_84:MULT_X_SUM_1;
signal  MULTS_1_85:MULT_X_SUM_1;
signal  MULTS_1_86:MULT_X_SUM_1;
signal  MULTS_1_87:MULT_X_SUM_1;
signal  MULTS_1_88:MULT_X_SUM_1;
signal  MULTS_1_89:MULT_X_SUM_1;
signal  MULTS_1_90:MULT_X_SUM_1;
signal  MULTS_1_91:MULT_X_SUM_1;
signal  MULTS_1_92:MULT_X_SUM_1;
signal  MULTS_1_93:MULT_X_SUM_1;
signal  MULTS_1_94:MULT_X_SUM_1;
signal  MULTS_1_95:MULT_X_SUM_1;
signal  MULTS_1_96:MULT_X_SUM_1;
signal  MULTS_1_97:MULT_X_SUM_1;
signal  MULTS_1_98:MULT_X_SUM_1;
signal  MULTS_1_99:MULT_X_SUM_1;
signal  MULTS_1_100:MULT_X_SUM_1;
signal  MULTS_1_101:MULT_X_SUM_1;
signal  MULTS_1_102:MULT_X_SUM_1;
signal  MULTS_1_103:MULT_X_SUM_1;
signal  MULTS_1_104:MULT_X_SUM_1;
signal  MULTS_1_105:MULT_X_SUM_1;
signal  MULTS_1_106:MULT_X_SUM_1;
signal  MULTS_1_107:MULT_X_SUM_1;
signal  MULTS_1_108:MULT_X_SUM_1;
signal  MULTS_1_109:MULT_X_SUM_1;
signal  MULTS_1_110:MULT_X_SUM_1;
signal  MULTS_1_111:MULT_X_SUM_1;
signal  MULTS_1_112:MULT_X_SUM_1;
signal  MULTS_1_113:MULT_X_SUM_1;
signal  MULTS_1_114:MULT_X_SUM_1;
signal  MULTS_1_115:MULT_X_SUM_1;
signal  MULTS_1_116:MULT_X_SUM_1;
signal  MULTS_1_117:MULT_X_SUM_1;
signal  MULTS_1_118:MULT_X_SUM_1;
signal  MULTS_1_119:MULT_X_SUM_1;
signal  MULTS_1_120:MULT_X_SUM_1;
type    MULT_X_SUM_2	is array (0 to FEATURE_MAPS-1) of signed(PRECISION-1 downto 0);
signal  EN_SUM_MULT_2	: std_logic;
signal  MULTS_2_1:MULT_X_SUM_2;
signal  MULTS_2_2:MULT_X_SUM_2;
signal  MULTS_2_3:MULT_X_SUM_2;
signal  MULTS_2_4:MULT_X_SUM_2;
signal  MULTS_2_5:MULT_X_SUM_2;
signal  MULTS_2_6:MULT_X_SUM_2;
signal  MULTS_2_7:MULT_X_SUM_2;
signal  MULTS_2_8:MULT_X_SUM_2;
signal  MULTS_2_9:MULT_X_SUM_2;
signal  MULTS_2_10:MULT_X_SUM_2;
signal  MULTS_2_11:MULT_X_SUM_2;
signal  MULTS_2_12:MULT_X_SUM_2;
signal  MULTS_2_13:MULT_X_SUM_2;
signal  MULTS_2_14:MULT_X_SUM_2;
signal  MULTS_2_15:MULT_X_SUM_2;
signal  MULTS_2_16:MULT_X_SUM_2;
signal  MULTS_2_17:MULT_X_SUM_2;
signal  MULTS_2_18:MULT_X_SUM_2;
signal  MULTS_2_19:MULT_X_SUM_2;
signal  MULTS_2_20:MULT_X_SUM_2;
signal  MULTS_2_21:MULT_X_SUM_2;
signal  MULTS_2_22:MULT_X_SUM_2;
signal  MULTS_2_23:MULT_X_SUM_2;
signal  MULTS_2_24:MULT_X_SUM_2;
signal  MULTS_2_25:MULT_X_SUM_2;
signal  MULTS_2_26:MULT_X_SUM_2;
signal  MULTS_2_27:MULT_X_SUM_2;
signal  MULTS_2_28:MULT_X_SUM_2;
signal  MULTS_2_29:MULT_X_SUM_2;
signal  MULTS_2_30:MULT_X_SUM_2;
signal  MULTS_2_31:MULT_X_SUM_2;
signal  MULTS_2_32:MULT_X_SUM_2;
signal  MULTS_2_33:MULT_X_SUM_2;
signal  MULTS_2_34:MULT_X_SUM_2;
signal  MULTS_2_35:MULT_X_SUM_2;
signal  MULTS_2_36:MULT_X_SUM_2;
signal  MULTS_2_37:MULT_X_SUM_2;
signal  MULTS_2_38:MULT_X_SUM_2;
signal  MULTS_2_39:MULT_X_SUM_2;
signal  MULTS_2_40:MULT_X_SUM_2;
signal  MULTS_2_41:MULT_X_SUM_2;
signal  MULTS_2_42:MULT_X_SUM_2;
signal  MULTS_2_43:MULT_X_SUM_2;
signal  MULTS_2_44:MULT_X_SUM_2;
signal  MULTS_2_45:MULT_X_SUM_2;
signal  MULTS_2_46:MULT_X_SUM_2;
signal  MULTS_2_47:MULT_X_SUM_2;
signal  MULTS_2_48:MULT_X_SUM_2;
signal  MULTS_2_49:MULT_X_SUM_2;
signal  MULTS_2_50:MULT_X_SUM_2;
signal  MULTS_2_51:MULT_X_SUM_2;
signal  MULTS_2_52:MULT_X_SUM_2;
signal  MULTS_2_53:MULT_X_SUM_2;
signal  MULTS_2_54:MULT_X_SUM_2;
signal  MULTS_2_55:MULT_X_SUM_2;
signal  MULTS_2_56:MULT_X_SUM_2;
signal  MULTS_2_57:MULT_X_SUM_2;
signal  MULTS_2_58:MULT_X_SUM_2;
signal  MULTS_2_59:MULT_X_SUM_2;
signal  MULTS_2_60:MULT_X_SUM_2;
signal  MULTS_2_61:MULT_X_SUM_2;
signal  MULTS_2_62:MULT_X_SUM_2;
signal  MULTS_2_63:MULT_X_SUM_2;
signal  MULTS_2_64:MULT_X_SUM_2;
signal  MULTS_2_65:MULT_X_SUM_2;
signal  MULTS_2_66:MULT_X_SUM_2;
signal  MULTS_2_67:MULT_X_SUM_2;
signal  MULTS_2_68:MULT_X_SUM_2;
signal  MULTS_2_69:MULT_X_SUM_2;
signal  MULTS_2_70:MULT_X_SUM_2;
signal  MULTS_2_71:MULT_X_SUM_2;
signal  MULTS_2_72:MULT_X_SUM_2;
signal  MULTS_2_73:MULT_X_SUM_2;
signal  MULTS_2_74:MULT_X_SUM_2;
signal  MULTS_2_75:MULT_X_SUM_2;
signal  MULTS_2_76:MULT_X_SUM_2;
signal  MULTS_2_77:MULT_X_SUM_2;
signal  MULTS_2_78:MULT_X_SUM_2;
signal  MULTS_2_79:MULT_X_SUM_2;
signal  MULTS_2_80:MULT_X_SUM_2;
signal  MULTS_2_81:MULT_X_SUM_2;
signal  MULTS_2_82:MULT_X_SUM_2;
signal  MULTS_2_83:MULT_X_SUM_2;
signal  MULTS_2_84:MULT_X_SUM_2;
signal  MULTS_2_85:MULT_X_SUM_2;
signal  MULTS_2_86:MULT_X_SUM_2;
signal  MULTS_2_87:MULT_X_SUM_2;
signal  MULTS_2_88:MULT_X_SUM_2;
signal  MULTS_2_89:MULT_X_SUM_2;
signal  MULTS_2_90:MULT_X_SUM_2;
signal  MULTS_2_91:MULT_X_SUM_2;
signal  MULTS_2_92:MULT_X_SUM_2;
signal  MULTS_2_93:MULT_X_SUM_2;
signal  MULTS_2_94:MULT_X_SUM_2;
signal  MULTS_2_95:MULT_X_SUM_2;
signal  MULTS_2_96:MULT_X_SUM_2;
signal  MULTS_2_97:MULT_X_SUM_2;
signal  MULTS_2_98:MULT_X_SUM_2;
signal  MULTS_2_99:MULT_X_SUM_2;
signal  MULTS_2_100:MULT_X_SUM_2;
signal  MULTS_2_101:MULT_X_SUM_2;
signal  MULTS_2_102:MULT_X_SUM_2;
signal  MULTS_2_103:MULT_X_SUM_2;
signal  MULTS_2_104:MULT_X_SUM_2;
signal  MULTS_2_105:MULT_X_SUM_2;
signal  MULTS_2_106:MULT_X_SUM_2;
signal  MULTS_2_107:MULT_X_SUM_2;
signal  MULTS_2_108:MULT_X_SUM_2;
signal  MULTS_2_109:MULT_X_SUM_2;
signal  MULTS_2_110:MULT_X_SUM_2;
signal  MULTS_2_111:MULT_X_SUM_2;
signal  MULTS_2_112:MULT_X_SUM_2;
signal  MULTS_2_113:MULT_X_SUM_2;
signal  MULTS_2_114:MULT_X_SUM_2;
signal  MULTS_2_115:MULT_X_SUM_2;
signal  MULTS_2_116:MULT_X_SUM_2;
signal  MULTS_2_117:MULT_X_SUM_2;
signal  MULTS_2_118:MULT_X_SUM_2;
signal  MULTS_2_119:MULT_X_SUM_2;
signal  MULTS_2_120:MULT_X_SUM_2;
type    MULT_X_SUM_3	is array (0 to FEATURE_MAPS-1) of signed(PRECISION-1 downto 0);
signal  EN_SUM_MULT_3	: std_logic;
signal  MULTS_3_1:MULT_X_SUM_3;
signal  MULTS_3_2:MULT_X_SUM_3;
signal  MULTS_3_3:MULT_X_SUM_3;
signal  MULTS_3_4:MULT_X_SUM_3;
signal  MULTS_3_5:MULT_X_SUM_3;
signal  MULTS_3_6:MULT_X_SUM_3;
signal  MULTS_3_7:MULT_X_SUM_3;
signal  MULTS_3_8:MULT_X_SUM_3;
signal  MULTS_3_9:MULT_X_SUM_3;
signal  MULTS_3_10:MULT_X_SUM_3;
signal  MULTS_3_11:MULT_X_SUM_3;
signal  MULTS_3_12:MULT_X_SUM_3;
signal  MULTS_3_13:MULT_X_SUM_3;
signal  MULTS_3_14:MULT_X_SUM_3;
signal  MULTS_3_15:MULT_X_SUM_3;
signal  MULTS_3_16:MULT_X_SUM_3;
signal  MULTS_3_17:MULT_X_SUM_3;
signal  MULTS_3_18:MULT_X_SUM_3;
signal  MULTS_3_19:MULT_X_SUM_3;
signal  MULTS_3_20:MULT_X_SUM_3;
signal  MULTS_3_21:MULT_X_SUM_3;
signal  MULTS_3_22:MULT_X_SUM_3;
signal  MULTS_3_23:MULT_X_SUM_3;
signal  MULTS_3_24:MULT_X_SUM_3;
signal  MULTS_3_25:MULT_X_SUM_3;
signal  MULTS_3_26:MULT_X_SUM_3;
signal  MULTS_3_27:MULT_X_SUM_3;
signal  MULTS_3_28:MULT_X_SUM_3;
signal  MULTS_3_29:MULT_X_SUM_3;
signal  MULTS_3_30:MULT_X_SUM_3;
signal  MULTS_3_31:MULT_X_SUM_3;
signal  MULTS_3_32:MULT_X_SUM_3;
signal  MULTS_3_33:MULT_X_SUM_3;
signal  MULTS_3_34:MULT_X_SUM_3;
signal  MULTS_3_35:MULT_X_SUM_3;
signal  MULTS_3_36:MULT_X_SUM_3;
signal  MULTS_3_37:MULT_X_SUM_3;
signal  MULTS_3_38:MULT_X_SUM_3;
signal  MULTS_3_39:MULT_X_SUM_3;
signal  MULTS_3_40:MULT_X_SUM_3;
signal  MULTS_3_41:MULT_X_SUM_3;
signal  MULTS_3_42:MULT_X_SUM_3;
signal  MULTS_3_43:MULT_X_SUM_3;
signal  MULTS_3_44:MULT_X_SUM_3;
signal  MULTS_3_45:MULT_X_SUM_3;
signal  MULTS_3_46:MULT_X_SUM_3;
signal  MULTS_3_47:MULT_X_SUM_3;
signal  MULTS_3_48:MULT_X_SUM_3;
signal  MULTS_3_49:MULT_X_SUM_3;
signal  MULTS_3_50:MULT_X_SUM_3;
signal  MULTS_3_51:MULT_X_SUM_3;
signal  MULTS_3_52:MULT_X_SUM_3;
signal  MULTS_3_53:MULT_X_SUM_3;
signal  MULTS_3_54:MULT_X_SUM_3;
signal  MULTS_3_55:MULT_X_SUM_3;
signal  MULTS_3_56:MULT_X_SUM_3;
signal  MULTS_3_57:MULT_X_SUM_3;
signal  MULTS_3_58:MULT_X_SUM_3;
signal  MULTS_3_59:MULT_X_SUM_3;
signal  MULTS_3_60:MULT_X_SUM_3;
signal  MULTS_3_61:MULT_X_SUM_3;
signal  MULTS_3_62:MULT_X_SUM_3;
signal  MULTS_3_63:MULT_X_SUM_3;
signal  MULTS_3_64:MULT_X_SUM_3;
signal  MULTS_3_65:MULT_X_SUM_3;
signal  MULTS_3_66:MULT_X_SUM_3;
signal  MULTS_3_67:MULT_X_SUM_3;
signal  MULTS_3_68:MULT_X_SUM_3;
signal  MULTS_3_69:MULT_X_SUM_3;
signal  MULTS_3_70:MULT_X_SUM_3;
signal  MULTS_3_71:MULT_X_SUM_3;
signal  MULTS_3_72:MULT_X_SUM_3;
signal  MULTS_3_73:MULT_X_SUM_3;
signal  MULTS_3_74:MULT_X_SUM_3;
signal  MULTS_3_75:MULT_X_SUM_3;
signal  MULTS_3_76:MULT_X_SUM_3;
signal  MULTS_3_77:MULT_X_SUM_3;
signal  MULTS_3_78:MULT_X_SUM_3;
signal  MULTS_3_79:MULT_X_SUM_3;
signal  MULTS_3_80:MULT_X_SUM_3;
signal  MULTS_3_81:MULT_X_SUM_3;
signal  MULTS_3_82:MULT_X_SUM_3;
signal  MULTS_3_83:MULT_X_SUM_3;
signal  MULTS_3_84:MULT_X_SUM_3;
signal  MULTS_3_85:MULT_X_SUM_3;
signal  MULTS_3_86:MULT_X_SUM_3;
signal  MULTS_3_87:MULT_X_SUM_3;
signal  MULTS_3_88:MULT_X_SUM_3;
signal  MULTS_3_89:MULT_X_SUM_3;
signal  MULTS_3_90:MULT_X_SUM_3;
signal  MULTS_3_91:MULT_X_SUM_3;
signal  MULTS_3_92:MULT_X_SUM_3;
signal  MULTS_3_93:MULT_X_SUM_3;
signal  MULTS_3_94:MULT_X_SUM_3;
signal  MULTS_3_95:MULT_X_SUM_3;
signal  MULTS_3_96:MULT_X_SUM_3;
signal  MULTS_3_97:MULT_X_SUM_3;
signal  MULTS_3_98:MULT_X_SUM_3;
signal  MULTS_3_99:MULT_X_SUM_3;
signal  MULTS_3_100:MULT_X_SUM_3;
signal  MULTS_3_101:MULT_X_SUM_3;
signal  MULTS_3_102:MULT_X_SUM_3;
signal  MULTS_3_103:MULT_X_SUM_3;
signal  MULTS_3_104:MULT_X_SUM_3;
signal  MULTS_3_105:MULT_X_SUM_3;
signal  MULTS_3_106:MULT_X_SUM_3;
signal  MULTS_3_107:MULT_X_SUM_3;
signal  MULTS_3_108:MULT_X_SUM_3;
signal  MULTS_3_109:MULT_X_SUM_3;
signal  MULTS_3_110:MULT_X_SUM_3;
signal  MULTS_3_111:MULT_X_SUM_3;
signal  MULTS_3_112:MULT_X_SUM_3;
signal  MULTS_3_113:MULT_X_SUM_3;
signal  MULTS_3_114:MULT_X_SUM_3;
signal  MULTS_3_115:MULT_X_SUM_3;
signal  MULTS_3_116:MULT_X_SUM_3;
signal  MULTS_3_117:MULT_X_SUM_3;
signal  MULTS_3_118:MULT_X_SUM_3;
signal  MULTS_3_119:MULT_X_SUM_3;
signal  MULTS_3_120:MULT_X_SUM_3;
type    MULT_X_SUM_4	is array (0 to FEATURE_MAPS-1) of signed(PRECISION-1 downto 0);
signal  EN_SUM_MULT_4	: std_logic;
signal  MULTS_4_1:MULT_X_SUM_4;
signal  MULTS_4_2:MULT_X_SUM_4;
signal  MULTS_4_3:MULT_X_SUM_4;
signal  MULTS_4_4:MULT_X_SUM_4;
signal  MULTS_4_5:MULT_X_SUM_4;
signal  MULTS_4_6:MULT_X_SUM_4;
signal  MULTS_4_7:MULT_X_SUM_4;
signal  MULTS_4_8:MULT_X_SUM_4;
signal  MULTS_4_9:MULT_X_SUM_4;
signal  MULTS_4_10:MULT_X_SUM_4;
signal  MULTS_4_11:MULT_X_SUM_4;
signal  MULTS_4_12:MULT_X_SUM_4;
signal  MULTS_4_13:MULT_X_SUM_4;
signal  MULTS_4_14:MULT_X_SUM_4;
signal  MULTS_4_15:MULT_X_SUM_4;
signal  MULTS_4_16:MULT_X_SUM_4;
signal  MULTS_4_17:MULT_X_SUM_4;
signal  MULTS_4_18:MULT_X_SUM_4;
signal  MULTS_4_19:MULT_X_SUM_4;
signal  MULTS_4_20:MULT_X_SUM_4;
signal  MULTS_4_21:MULT_X_SUM_4;
signal  MULTS_4_22:MULT_X_SUM_4;
signal  MULTS_4_23:MULT_X_SUM_4;
signal  MULTS_4_24:MULT_X_SUM_4;
signal  MULTS_4_25:MULT_X_SUM_4;
signal  MULTS_4_26:MULT_X_SUM_4;
signal  MULTS_4_27:MULT_X_SUM_4;
signal  MULTS_4_28:MULT_X_SUM_4;
signal  MULTS_4_29:MULT_X_SUM_4;
signal  MULTS_4_30:MULT_X_SUM_4;
signal  MULTS_4_31:MULT_X_SUM_4;
signal  MULTS_4_32:MULT_X_SUM_4;
signal  MULTS_4_33:MULT_X_SUM_4;
signal  MULTS_4_34:MULT_X_SUM_4;
signal  MULTS_4_35:MULT_X_SUM_4;
signal  MULTS_4_36:MULT_X_SUM_4;
signal  MULTS_4_37:MULT_X_SUM_4;
signal  MULTS_4_38:MULT_X_SUM_4;
signal  MULTS_4_39:MULT_X_SUM_4;
signal  MULTS_4_40:MULT_X_SUM_4;
signal  MULTS_4_41:MULT_X_SUM_4;
signal  MULTS_4_42:MULT_X_SUM_4;
signal  MULTS_4_43:MULT_X_SUM_4;
signal  MULTS_4_44:MULT_X_SUM_4;
signal  MULTS_4_45:MULT_X_SUM_4;
signal  MULTS_4_46:MULT_X_SUM_4;
signal  MULTS_4_47:MULT_X_SUM_4;
signal  MULTS_4_48:MULT_X_SUM_4;
signal  MULTS_4_49:MULT_X_SUM_4;
signal  MULTS_4_50:MULT_X_SUM_4;
signal  MULTS_4_51:MULT_X_SUM_4;
signal  MULTS_4_52:MULT_X_SUM_4;
signal  MULTS_4_53:MULT_X_SUM_4;
signal  MULTS_4_54:MULT_X_SUM_4;
signal  MULTS_4_55:MULT_X_SUM_4;
signal  MULTS_4_56:MULT_X_SUM_4;
signal  MULTS_4_57:MULT_X_SUM_4;
signal  MULTS_4_58:MULT_X_SUM_4;
signal  MULTS_4_59:MULT_X_SUM_4;
signal  MULTS_4_60:MULT_X_SUM_4;
signal  MULTS_4_61:MULT_X_SUM_4;
signal  MULTS_4_62:MULT_X_SUM_4;
signal  MULTS_4_63:MULT_X_SUM_4;
signal  MULTS_4_64:MULT_X_SUM_4;
signal  MULTS_4_65:MULT_X_SUM_4;
signal  MULTS_4_66:MULT_X_SUM_4;
signal  MULTS_4_67:MULT_X_SUM_4;
signal  MULTS_4_68:MULT_X_SUM_4;
signal  MULTS_4_69:MULT_X_SUM_4;
signal  MULTS_4_70:MULT_X_SUM_4;
signal  MULTS_4_71:MULT_X_SUM_4;
signal  MULTS_4_72:MULT_X_SUM_4;
signal  MULTS_4_73:MULT_X_SUM_4;
signal  MULTS_4_74:MULT_X_SUM_4;
signal  MULTS_4_75:MULT_X_SUM_4;
signal  MULTS_4_76:MULT_X_SUM_4;
signal  MULTS_4_77:MULT_X_SUM_4;
signal  MULTS_4_78:MULT_X_SUM_4;
signal  MULTS_4_79:MULT_X_SUM_4;
signal  MULTS_4_80:MULT_X_SUM_4;
signal  MULTS_4_81:MULT_X_SUM_4;
signal  MULTS_4_82:MULT_X_SUM_4;
signal  MULTS_4_83:MULT_X_SUM_4;
signal  MULTS_4_84:MULT_X_SUM_4;
signal  MULTS_4_85:MULT_X_SUM_4;
signal  MULTS_4_86:MULT_X_SUM_4;
signal  MULTS_4_87:MULT_X_SUM_4;
signal  MULTS_4_88:MULT_X_SUM_4;
signal  MULTS_4_89:MULT_X_SUM_4;
signal  MULTS_4_90:MULT_X_SUM_4;
signal  MULTS_4_91:MULT_X_SUM_4;
signal  MULTS_4_92:MULT_X_SUM_4;
signal  MULTS_4_93:MULT_X_SUM_4;
signal  MULTS_4_94:MULT_X_SUM_4;
signal  MULTS_4_95:MULT_X_SUM_4;
signal  MULTS_4_96:MULT_X_SUM_4;
signal  MULTS_4_97:MULT_X_SUM_4;
signal  MULTS_4_98:MULT_X_SUM_4;
signal  MULTS_4_99:MULT_X_SUM_4;
signal  MULTS_4_100:MULT_X_SUM_4;
signal  MULTS_4_101:MULT_X_SUM_4;
signal  MULTS_4_102:MULT_X_SUM_4;
signal  MULTS_4_103:MULT_X_SUM_4;
signal  MULTS_4_104:MULT_X_SUM_4;
signal  MULTS_4_105:MULT_X_SUM_4;
signal  MULTS_4_106:MULT_X_SUM_4;
signal  MULTS_4_107:MULT_X_SUM_4;
signal  MULTS_4_108:MULT_X_SUM_4;
signal  MULTS_4_109:MULT_X_SUM_4;
signal  MULTS_4_110:MULT_X_SUM_4;
signal  MULTS_4_111:MULT_X_SUM_4;
signal  MULTS_4_112:MULT_X_SUM_4;
signal  MULTS_4_113:MULT_X_SUM_4;
signal  MULTS_4_114:MULT_X_SUM_4;
signal  MULTS_4_115:MULT_X_SUM_4;
signal  MULTS_4_116:MULT_X_SUM_4;
signal  MULTS_4_117:MULT_X_SUM_4;
signal  MULTS_4_118:MULT_X_SUM_4;
signal  MULTS_4_119:MULT_X_SUM_4;
signal  MULTS_4_120:MULT_X_SUM_4;
type    MULT_X_SUM_5	is array (0 to FEATURE_MAPS-1) of signed(PRECISION-1 downto 0);
signal  EN_SUM_MULT_5	: std_logic;
signal  MULTS_5_1:MULT_X_SUM_5;
signal  MULTS_5_2:MULT_X_SUM_5;
signal  MULTS_5_3:MULT_X_SUM_5;
signal  MULTS_5_4:MULT_X_SUM_5;
signal  MULTS_5_5:MULT_X_SUM_5;
signal  MULTS_5_6:MULT_X_SUM_5;
signal  MULTS_5_7:MULT_X_SUM_5;
signal  MULTS_5_8:MULT_X_SUM_5;
signal  MULTS_5_9:MULT_X_SUM_5;
signal  MULTS_5_10:MULT_X_SUM_5;
signal  MULTS_5_11:MULT_X_SUM_5;
signal  MULTS_5_12:MULT_X_SUM_5;
signal  MULTS_5_13:MULT_X_SUM_5;
signal  MULTS_5_14:MULT_X_SUM_5;
signal  MULTS_5_15:MULT_X_SUM_5;
signal  MULTS_5_16:MULT_X_SUM_5;
signal  MULTS_5_17:MULT_X_SUM_5;
signal  MULTS_5_18:MULT_X_SUM_5;
signal  MULTS_5_19:MULT_X_SUM_5;
signal  MULTS_5_20:MULT_X_SUM_5;
signal  MULTS_5_21:MULT_X_SUM_5;
signal  MULTS_5_22:MULT_X_SUM_5;
signal  MULTS_5_23:MULT_X_SUM_5;
signal  MULTS_5_24:MULT_X_SUM_5;
signal  MULTS_5_25:MULT_X_SUM_5;
signal  MULTS_5_26:MULT_X_SUM_5;
signal  MULTS_5_27:MULT_X_SUM_5;
signal  MULTS_5_28:MULT_X_SUM_5;
signal  MULTS_5_29:MULT_X_SUM_5;
signal  MULTS_5_30:MULT_X_SUM_5;
signal  MULTS_5_31:MULT_X_SUM_5;
signal  MULTS_5_32:MULT_X_SUM_5;
signal  MULTS_5_33:MULT_X_SUM_5;
signal  MULTS_5_34:MULT_X_SUM_5;
signal  MULTS_5_35:MULT_X_SUM_5;
signal  MULTS_5_36:MULT_X_SUM_5;
signal  MULTS_5_37:MULT_X_SUM_5;
signal  MULTS_5_38:MULT_X_SUM_5;
signal  MULTS_5_39:MULT_X_SUM_5;
signal  MULTS_5_40:MULT_X_SUM_5;
signal  MULTS_5_41:MULT_X_SUM_5;
signal  MULTS_5_42:MULT_X_SUM_5;
signal  MULTS_5_43:MULT_X_SUM_5;
signal  MULTS_5_44:MULT_X_SUM_5;
signal  MULTS_5_45:MULT_X_SUM_5;
signal  MULTS_5_46:MULT_X_SUM_5;
signal  MULTS_5_47:MULT_X_SUM_5;
signal  MULTS_5_48:MULT_X_SUM_5;
signal  MULTS_5_49:MULT_X_SUM_5;
signal  MULTS_5_50:MULT_X_SUM_5;
signal  MULTS_5_51:MULT_X_SUM_5;
signal  MULTS_5_52:MULT_X_SUM_5;
signal  MULTS_5_53:MULT_X_SUM_5;
signal  MULTS_5_54:MULT_X_SUM_5;
signal  MULTS_5_55:MULT_X_SUM_5;
signal  MULTS_5_56:MULT_X_SUM_5;
signal  MULTS_5_57:MULT_X_SUM_5;
signal  MULTS_5_58:MULT_X_SUM_5;
signal  MULTS_5_59:MULT_X_SUM_5;
signal  MULTS_5_60:MULT_X_SUM_5;
signal  MULTS_5_61:MULT_X_SUM_5;
signal  MULTS_5_62:MULT_X_SUM_5;
signal  MULTS_5_63:MULT_X_SUM_5;
signal  MULTS_5_64:MULT_X_SUM_5;
signal  MULTS_5_65:MULT_X_SUM_5;
signal  MULTS_5_66:MULT_X_SUM_5;
signal  MULTS_5_67:MULT_X_SUM_5;
signal  MULTS_5_68:MULT_X_SUM_5;
signal  MULTS_5_69:MULT_X_SUM_5;
signal  MULTS_5_70:MULT_X_SUM_5;
signal  MULTS_5_71:MULT_X_SUM_5;
signal  MULTS_5_72:MULT_X_SUM_5;
signal  MULTS_5_73:MULT_X_SUM_5;
signal  MULTS_5_74:MULT_X_SUM_5;
signal  MULTS_5_75:MULT_X_SUM_5;
signal  MULTS_5_76:MULT_X_SUM_5;
signal  MULTS_5_77:MULT_X_SUM_5;
signal  MULTS_5_78:MULT_X_SUM_5;
signal  MULTS_5_79:MULT_X_SUM_5;
signal  MULTS_5_80:MULT_X_SUM_5;
signal  MULTS_5_81:MULT_X_SUM_5;
signal  MULTS_5_82:MULT_X_SUM_5;
signal  MULTS_5_83:MULT_X_SUM_5;
signal  MULTS_5_84:MULT_X_SUM_5;
signal  MULTS_5_85:MULT_X_SUM_5;
signal  MULTS_5_86:MULT_X_SUM_5;
signal  MULTS_5_87:MULT_X_SUM_5;
signal  MULTS_5_88:MULT_X_SUM_5;
signal  MULTS_5_89:MULT_X_SUM_5;
signal  MULTS_5_90:MULT_X_SUM_5;
signal  MULTS_5_91:MULT_X_SUM_5;
signal  MULTS_5_92:MULT_X_SUM_5;
signal  MULTS_5_93:MULT_X_SUM_5;
signal  MULTS_5_94:MULT_X_SUM_5;
signal  MULTS_5_95:MULT_X_SUM_5;
signal  MULTS_5_96:MULT_X_SUM_5;
signal  MULTS_5_97:MULT_X_SUM_5;
signal  MULTS_5_98:MULT_X_SUM_5;
signal  MULTS_5_99:MULT_X_SUM_5;
signal  MULTS_5_100:MULT_X_SUM_5;
signal  MULTS_5_101:MULT_X_SUM_5;
signal  MULTS_5_102:MULT_X_SUM_5;
signal  MULTS_5_103:MULT_X_SUM_5;
signal  MULTS_5_104:MULT_X_SUM_5;
signal  MULTS_5_105:MULT_X_SUM_5;
signal  MULTS_5_106:MULT_X_SUM_5;
signal  MULTS_5_107:MULT_X_SUM_5;
signal  MULTS_5_108:MULT_X_SUM_5;
signal  MULTS_5_109:MULT_X_SUM_5;
signal  MULTS_5_110:MULT_X_SUM_5;
signal  MULTS_5_111:MULT_X_SUM_5;
signal  MULTS_5_112:MULT_X_SUM_5;
signal  MULTS_5_113:MULT_X_SUM_5;
signal  MULTS_5_114:MULT_X_SUM_5;
signal  MULTS_5_115:MULT_X_SUM_5;
signal  MULTS_5_116:MULT_X_SUM_5;
signal  MULTS_5_117:MULT_X_SUM_5;
signal  MULTS_5_118:MULT_X_SUM_5;
signal  MULTS_5_119:MULT_X_SUM_5;
signal  MULTS_5_120:MULT_X_SUM_5;
type    MULT_X_SUM_6	is array (0 to FEATURE_MAPS-1) of signed(PRECISION-1 downto 0);
signal  EN_SUM_MULT_6	: std_logic;
signal  MULTS_6_1:MULT_X_SUM_6;
signal  MULTS_6_2:MULT_X_SUM_6;
signal  MULTS_6_3:MULT_X_SUM_6;
signal  MULTS_6_4:MULT_X_SUM_6;
signal  MULTS_6_5:MULT_X_SUM_6;
signal  MULTS_6_6:MULT_X_SUM_6;
signal  MULTS_6_7:MULT_X_SUM_6;
signal  MULTS_6_8:MULT_X_SUM_6;
signal  MULTS_6_9:MULT_X_SUM_6;
signal  MULTS_6_10:MULT_X_SUM_6;
signal  MULTS_6_11:MULT_X_SUM_6;
signal  MULTS_6_12:MULT_X_SUM_6;
signal  MULTS_6_13:MULT_X_SUM_6;
signal  MULTS_6_14:MULT_X_SUM_6;
signal  MULTS_6_15:MULT_X_SUM_6;
signal  MULTS_6_16:MULT_X_SUM_6;
signal  MULTS_6_17:MULT_X_SUM_6;
signal  MULTS_6_18:MULT_X_SUM_6;
signal  MULTS_6_19:MULT_X_SUM_6;
signal  MULTS_6_20:MULT_X_SUM_6;
signal  MULTS_6_21:MULT_X_SUM_6;
signal  MULTS_6_22:MULT_X_SUM_6;
signal  MULTS_6_23:MULT_X_SUM_6;
signal  MULTS_6_24:MULT_X_SUM_6;
signal  MULTS_6_25:MULT_X_SUM_6;
signal  MULTS_6_26:MULT_X_SUM_6;
signal  MULTS_6_27:MULT_X_SUM_6;
signal  MULTS_6_28:MULT_X_SUM_6;
signal  MULTS_6_29:MULT_X_SUM_6;
signal  MULTS_6_30:MULT_X_SUM_6;
signal  MULTS_6_31:MULT_X_SUM_6;
signal  MULTS_6_32:MULT_X_SUM_6;
signal  MULTS_6_33:MULT_X_SUM_6;
signal  MULTS_6_34:MULT_X_SUM_6;
signal  MULTS_6_35:MULT_X_SUM_6;
signal  MULTS_6_36:MULT_X_SUM_6;
signal  MULTS_6_37:MULT_X_SUM_6;
signal  MULTS_6_38:MULT_X_SUM_6;
signal  MULTS_6_39:MULT_X_SUM_6;
signal  MULTS_6_40:MULT_X_SUM_6;
signal  MULTS_6_41:MULT_X_SUM_6;
signal  MULTS_6_42:MULT_X_SUM_6;
signal  MULTS_6_43:MULT_X_SUM_6;
signal  MULTS_6_44:MULT_X_SUM_6;
signal  MULTS_6_45:MULT_X_SUM_6;
signal  MULTS_6_46:MULT_X_SUM_6;
signal  MULTS_6_47:MULT_X_SUM_6;
signal  MULTS_6_48:MULT_X_SUM_6;
signal  MULTS_6_49:MULT_X_SUM_6;
signal  MULTS_6_50:MULT_X_SUM_6;
signal  MULTS_6_51:MULT_X_SUM_6;
signal  MULTS_6_52:MULT_X_SUM_6;
signal  MULTS_6_53:MULT_X_SUM_6;
signal  MULTS_6_54:MULT_X_SUM_6;
signal  MULTS_6_55:MULT_X_SUM_6;
signal  MULTS_6_56:MULT_X_SUM_6;
signal  MULTS_6_57:MULT_X_SUM_6;
signal  MULTS_6_58:MULT_X_SUM_6;
signal  MULTS_6_59:MULT_X_SUM_6;
signal  MULTS_6_60:MULT_X_SUM_6;
signal  MULTS_6_61:MULT_X_SUM_6;
signal  MULTS_6_62:MULT_X_SUM_6;
signal  MULTS_6_63:MULT_X_SUM_6;
signal  MULTS_6_64:MULT_X_SUM_6;
signal  MULTS_6_65:MULT_X_SUM_6;
signal  MULTS_6_66:MULT_X_SUM_6;
signal  MULTS_6_67:MULT_X_SUM_6;
signal  MULTS_6_68:MULT_X_SUM_6;
signal  MULTS_6_69:MULT_X_SUM_6;
signal  MULTS_6_70:MULT_X_SUM_6;
signal  MULTS_6_71:MULT_X_SUM_6;
signal  MULTS_6_72:MULT_X_SUM_6;
signal  MULTS_6_73:MULT_X_SUM_6;
signal  MULTS_6_74:MULT_X_SUM_6;
signal  MULTS_6_75:MULT_X_SUM_6;
signal  MULTS_6_76:MULT_X_SUM_6;
signal  MULTS_6_77:MULT_X_SUM_6;
signal  MULTS_6_78:MULT_X_SUM_6;
signal  MULTS_6_79:MULT_X_SUM_6;
signal  MULTS_6_80:MULT_X_SUM_6;
signal  MULTS_6_81:MULT_X_SUM_6;
signal  MULTS_6_82:MULT_X_SUM_6;
signal  MULTS_6_83:MULT_X_SUM_6;
signal  MULTS_6_84:MULT_X_SUM_6;
signal  MULTS_6_85:MULT_X_SUM_6;
signal  MULTS_6_86:MULT_X_SUM_6;
signal  MULTS_6_87:MULT_X_SUM_6;
signal  MULTS_6_88:MULT_X_SUM_6;
signal  MULTS_6_89:MULT_X_SUM_6;
signal  MULTS_6_90:MULT_X_SUM_6;
signal  MULTS_6_91:MULT_X_SUM_6;
signal  MULTS_6_92:MULT_X_SUM_6;
signal  MULTS_6_93:MULT_X_SUM_6;
signal  MULTS_6_94:MULT_X_SUM_6;
signal  MULTS_6_95:MULT_X_SUM_6;
signal  MULTS_6_96:MULT_X_SUM_6;
signal  MULTS_6_97:MULT_X_SUM_6;
signal  MULTS_6_98:MULT_X_SUM_6;
signal  MULTS_6_99:MULT_X_SUM_6;
signal  MULTS_6_100:MULT_X_SUM_6;
signal  MULTS_6_101:MULT_X_SUM_6;
signal  MULTS_6_102:MULT_X_SUM_6;
signal  MULTS_6_103:MULT_X_SUM_6;
signal  MULTS_6_104:MULT_X_SUM_6;
signal  MULTS_6_105:MULT_X_SUM_6;
signal  MULTS_6_106:MULT_X_SUM_6;
signal  MULTS_6_107:MULT_X_SUM_6;
signal  MULTS_6_108:MULT_X_SUM_6;
signal  MULTS_6_109:MULT_X_SUM_6;
signal  MULTS_6_110:MULT_X_SUM_6;
signal  MULTS_6_111:MULT_X_SUM_6;
signal  MULTS_6_112:MULT_X_SUM_6;
signal  MULTS_6_113:MULT_X_SUM_6;
signal  MULTS_6_114:MULT_X_SUM_6;
signal  MULTS_6_115:MULT_X_SUM_6;
signal  MULTS_6_116:MULT_X_SUM_6;
signal  MULTS_6_117:MULT_X_SUM_6;
signal  MULTS_6_118:MULT_X_SUM_6;
signal  MULTS_6_119:MULT_X_SUM_6;
signal  MULTS_6_120:MULT_X_SUM_6;
type    MULT_X_SUM_7	is array (0 to FEATURE_MAPS-1) of signed(PRECISION-1 downto 0);
signal  EN_SUM_MULT_7	: std_logic;
signal  MULTS_7_1:MULT_X_SUM_7;
signal  MULTS_7_2:MULT_X_SUM_7;
signal  MULTS_7_3:MULT_X_SUM_7;
signal  MULTS_7_4:MULT_X_SUM_7;
signal  MULTS_7_5:MULT_X_SUM_7;
signal  MULTS_7_6:MULT_X_SUM_7;
signal  MULTS_7_7:MULT_X_SUM_7;
signal  MULTS_7_8:MULT_X_SUM_7;
signal  MULTS_7_9:MULT_X_SUM_7;
signal  MULTS_7_10:MULT_X_SUM_7;
signal  MULTS_7_11:MULT_X_SUM_7;
signal  MULTS_7_12:MULT_X_SUM_7;
signal  MULTS_7_13:MULT_X_SUM_7;
signal  MULTS_7_14:MULT_X_SUM_7;
signal  MULTS_7_15:MULT_X_SUM_7;
signal  MULTS_7_16:MULT_X_SUM_7;
signal  MULTS_7_17:MULT_X_SUM_7;
signal  MULTS_7_18:MULT_X_SUM_7;
signal  MULTS_7_19:MULT_X_SUM_7;
signal  MULTS_7_20:MULT_X_SUM_7;
signal  MULTS_7_21:MULT_X_SUM_7;
signal  MULTS_7_22:MULT_X_SUM_7;
signal  MULTS_7_23:MULT_X_SUM_7;
signal  MULTS_7_24:MULT_X_SUM_7;
signal  MULTS_7_25:MULT_X_SUM_7;
signal  MULTS_7_26:MULT_X_SUM_7;
signal  MULTS_7_27:MULT_X_SUM_7;
signal  MULTS_7_28:MULT_X_SUM_7;
signal  MULTS_7_29:MULT_X_SUM_7;
signal  MULTS_7_30:MULT_X_SUM_7;
signal  MULTS_7_31:MULT_X_SUM_7;
signal  MULTS_7_32:MULT_X_SUM_7;
signal  MULTS_7_33:MULT_X_SUM_7;
signal  MULTS_7_34:MULT_X_SUM_7;
signal  MULTS_7_35:MULT_X_SUM_7;
signal  MULTS_7_36:MULT_X_SUM_7;
signal  MULTS_7_37:MULT_X_SUM_7;
signal  MULTS_7_38:MULT_X_SUM_7;
signal  MULTS_7_39:MULT_X_SUM_7;
signal  MULTS_7_40:MULT_X_SUM_7;
signal  MULTS_7_41:MULT_X_SUM_7;
signal  MULTS_7_42:MULT_X_SUM_7;
signal  MULTS_7_43:MULT_X_SUM_7;
signal  MULTS_7_44:MULT_X_SUM_7;
signal  MULTS_7_45:MULT_X_SUM_7;
signal  MULTS_7_46:MULT_X_SUM_7;
signal  MULTS_7_47:MULT_X_SUM_7;
signal  MULTS_7_48:MULT_X_SUM_7;
signal  MULTS_7_49:MULT_X_SUM_7;
signal  MULTS_7_50:MULT_X_SUM_7;
signal  MULTS_7_51:MULT_X_SUM_7;
signal  MULTS_7_52:MULT_X_SUM_7;
signal  MULTS_7_53:MULT_X_SUM_7;
signal  MULTS_7_54:MULT_X_SUM_7;
signal  MULTS_7_55:MULT_X_SUM_7;
signal  MULTS_7_56:MULT_X_SUM_7;
signal  MULTS_7_57:MULT_X_SUM_7;
signal  MULTS_7_58:MULT_X_SUM_7;
signal  MULTS_7_59:MULT_X_SUM_7;
signal  MULTS_7_60:MULT_X_SUM_7;
signal  MULTS_7_61:MULT_X_SUM_7;
signal  MULTS_7_62:MULT_X_SUM_7;
signal  MULTS_7_63:MULT_X_SUM_7;
signal  MULTS_7_64:MULT_X_SUM_7;
signal  MULTS_7_65:MULT_X_SUM_7;
signal  MULTS_7_66:MULT_X_SUM_7;
signal  MULTS_7_67:MULT_X_SUM_7;
signal  MULTS_7_68:MULT_X_SUM_7;
signal  MULTS_7_69:MULT_X_SUM_7;
signal  MULTS_7_70:MULT_X_SUM_7;
signal  MULTS_7_71:MULT_X_SUM_7;
signal  MULTS_7_72:MULT_X_SUM_7;
signal  MULTS_7_73:MULT_X_SUM_7;
signal  MULTS_7_74:MULT_X_SUM_7;
signal  MULTS_7_75:MULT_X_SUM_7;
signal  MULTS_7_76:MULT_X_SUM_7;
signal  MULTS_7_77:MULT_X_SUM_7;
signal  MULTS_7_78:MULT_X_SUM_7;
signal  MULTS_7_79:MULT_X_SUM_7;
signal  MULTS_7_80:MULT_X_SUM_7;
signal  MULTS_7_81:MULT_X_SUM_7;
signal  MULTS_7_82:MULT_X_SUM_7;
signal  MULTS_7_83:MULT_X_SUM_7;
signal  MULTS_7_84:MULT_X_SUM_7;
signal  MULTS_7_85:MULT_X_SUM_7;
signal  MULTS_7_86:MULT_X_SUM_7;
signal  MULTS_7_87:MULT_X_SUM_7;
signal  MULTS_7_88:MULT_X_SUM_7;
signal  MULTS_7_89:MULT_X_SUM_7;
signal  MULTS_7_90:MULT_X_SUM_7;
signal  MULTS_7_91:MULT_X_SUM_7;
signal  MULTS_7_92:MULT_X_SUM_7;
signal  MULTS_7_93:MULT_X_SUM_7;
signal  MULTS_7_94:MULT_X_SUM_7;
signal  MULTS_7_95:MULT_X_SUM_7;
signal  MULTS_7_96:MULT_X_SUM_7;
signal  MULTS_7_97:MULT_X_SUM_7;
signal  MULTS_7_98:MULT_X_SUM_7;
signal  MULTS_7_99:MULT_X_SUM_7;
signal  MULTS_7_100:MULT_X_SUM_7;
signal  MULTS_7_101:MULT_X_SUM_7;
signal  MULTS_7_102:MULT_X_SUM_7;
signal  MULTS_7_103:MULT_X_SUM_7;
signal  MULTS_7_104:MULT_X_SUM_7;
signal  MULTS_7_105:MULT_X_SUM_7;
signal  MULTS_7_106:MULT_X_SUM_7;
signal  MULTS_7_107:MULT_X_SUM_7;
signal  MULTS_7_108:MULT_X_SUM_7;
signal  MULTS_7_109:MULT_X_SUM_7;
signal  MULTS_7_110:MULT_X_SUM_7;
signal  MULTS_7_111:MULT_X_SUM_7;
signal  MULTS_7_112:MULT_X_SUM_7;
signal  MULTS_7_113:MULT_X_SUM_7;
signal  MULTS_7_114:MULT_X_SUM_7;
signal  MULTS_7_115:MULT_X_SUM_7;
signal  MULTS_7_116:MULT_X_SUM_7;
signal  MULTS_7_117:MULT_X_SUM_7;
signal  MULTS_7_118:MULT_X_SUM_7;
signal  MULTS_7_119:MULT_X_SUM_7;
signal  MULTS_7_120:MULT_X_SUM_7;



--------------------------------------------- FILTER HARDCODED CONSTANTS -WEIGHTS START--------------------------------

constant FMAP_1_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_1_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_2_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_3_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_4_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_5_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_6_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_7_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_8_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_9_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_1: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_2: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_3: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_4: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_5: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_6: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_7: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_8: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_9: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_10: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_11: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_12: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_13: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_14: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_15: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_16: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_17: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_18: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_19: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_20: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_21: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_22: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_23: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_24: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_25: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_26: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_27: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_28: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_29: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_30: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_31: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_32: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_33: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_34: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_35: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_36: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_37: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_38: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_39: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_40: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_41: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_42: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_43: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_44: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_45: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_46: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_47: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_48: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_49: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_50: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_51: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_52: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_53: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_54: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_55: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_56: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_57: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_58: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_59: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_60: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_61: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_62: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_63: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_64: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_65: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_66: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_67: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_68: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_69: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_70: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_71: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_72: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_73: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_74: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_75: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_76: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_77: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_78: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_79: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_80: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_81: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_82: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_83: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_84: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_85: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_86: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_87: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_88: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_89: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_90: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_91: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_92: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_93: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_94: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_95: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_96: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_97: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_98: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_99: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_100: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_101: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_102: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_103: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_104: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_105: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_106: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_107: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_108: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_109: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_110: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_111: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_112: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_113: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_114: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_115: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_116: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_117: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_118: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_119: signed(WEIGHT_SIZE- 1 downto 0):= "00001";
constant FMAP_10_120: signed(WEIGHT_SIZE- 1 downto 0):= "00001";

constant BIAS_VAL_1: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_2: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_3: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_4: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_5: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_6: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_7: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_8: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_9: signed (BIASES_SIZE-1 downto 0):="01";
constant BIAS_VAL_10: signed (BIASES_SIZE-1 downto 0):="01";


BEGIN
-------------------------------------------------------- ARCHITECTURE BEGIN--------------------------------------------------------

LAYER_7: process(CLK)


begin
------------------------------------------------ RESET AND PROCESS TOP START ------------------------------------------------------
if rising_edge(CLK) then
  if RST = '1' then
	-------------------FIXED SIGNALS RESET------------------------
    PIXEL_COUNT<=0;VALID_NXTLYR_PIX<=0;OUT_PIXEL_COUNT<=0;
    EN_NXT_LYR_7<='0';FRST_TIM_EN_7<='0';INTERNAL_RST<='0';
    Enable_MULT<='0';Enable_ADDER<='0';Enable_ReLU<='0';Enable_BIAS<='0';
    PADDING_count<=0;ROW_COUNT<=0;SIG_STRIDE<=STRIDE;COUNT_PIX<=0;

-------------------DYNAMIC SIGNALS RESET------------------------
    DOUT_BUF_1_7<=(others => '0');BIAS_1<=(others => '0');ReLU_1<=(others => '0');
    DOUT_BUF_2_7<=(others => '0');BIAS_2<=(others => '0');ReLU_2<=(others => '0');
    DOUT_BUF_3_7<=(others => '0');BIAS_3<=(others => '0');ReLU_3<=(others => '0');
    DOUT_BUF_4_7<=(others => '0');BIAS_4<=(others => '0');ReLU_4<=(others => '0');
    DOUT_BUF_5_7<=(others => '0');BIAS_5<=(others => '0');ReLU_5<=(others => '0');
    DOUT_BUF_6_7<=(others => '0');BIAS_6<=(others => '0');ReLU_6<=(others => '0');
    DOUT_BUF_7_7<=(others => '0');BIAS_7<=(others => '0');ReLU_7<=(others => '0');
    DOUT_BUF_8_7<=(others => '0');BIAS_8<=(others => '0');ReLU_8<=(others => '0');
    DOUT_BUF_9_7<=(others => '0');BIAS_9<=(others => '0');ReLU_9<=(others => '0');
    DOUT_BUF_10_7<=(others => '0');BIAS_10<=(others => '0');ReLU_10<=(others => '0');

    SUM_PIXELS_1<=(others=>'0');MULT_1<=((others=> (others=>'0')));
    SUM_PIXELS_2<=(others=>'0');MULT_2<=((others=> (others=>'0')));
    SUM_PIXELS_3<=(others=>'0');MULT_3<=((others=> (others=>'0')));
    SUM_PIXELS_4<=(others=>'0');MULT_4<=((others=> (others=>'0')));
    SUM_PIXELS_5<=(others=>'0');MULT_5<=((others=> (others=>'0')));
    SUM_PIXELS_6<=(others=>'0');MULT_6<=((others=> (others=>'0')));
    SUM_PIXELS_7<=(others=>'0');MULT_7<=((others=> (others=>'0')));
    SUM_PIXELS_8<=(others=>'0');MULT_8<=((others=> (others=>'0')));
    SUM_PIXELS_9<=(others=>'0');MULT_9<=((others=> (others=>'0')));
    SUM_PIXELS_10<=(others=>'0');MULT_10<=((others=> (others=>'0')));
    SUM_PIXELS_11<=(others=>'0');MULT_11<=((others=> (others=>'0')));
    SUM_PIXELS_12<=(others=>'0');MULT_12<=((others=> (others=>'0')));
    SUM_PIXELS_13<=(others=>'0');MULT_13<=((others=> (others=>'0')));
    SUM_PIXELS_14<=(others=>'0');MULT_14<=((others=> (others=>'0')));
    SUM_PIXELS_15<=(others=>'0');MULT_15<=((others=> (others=>'0')));
    SUM_PIXELS_16<=(others=>'0');MULT_16<=((others=> (others=>'0')));
    SUM_PIXELS_17<=(others=>'0');MULT_17<=((others=> (others=>'0')));
    SUM_PIXELS_18<=(others=>'0');MULT_18<=((others=> (others=>'0')));
    SUM_PIXELS_19<=(others=>'0');MULT_19<=((others=> (others=>'0')));
    SUM_PIXELS_20<=(others=>'0');MULT_20<=((others=> (others=>'0')));
    SUM_PIXELS_21<=(others=>'0');MULT_21<=((others=> (others=>'0')));
    SUM_PIXELS_22<=(others=>'0');MULT_22<=((others=> (others=>'0')));
    SUM_PIXELS_23<=(others=>'0');MULT_23<=((others=> (others=>'0')));
    SUM_PIXELS_24<=(others=>'0');MULT_24<=((others=> (others=>'0')));
    SUM_PIXELS_25<=(others=>'0');MULT_25<=((others=> (others=>'0')));
    SUM_PIXELS_26<=(others=>'0');MULT_26<=((others=> (others=>'0')));
    SUM_PIXELS_27<=(others=>'0');MULT_27<=((others=> (others=>'0')));
    SUM_PIXELS_28<=(others=>'0');MULT_28<=((others=> (others=>'0')));
    SUM_PIXELS_29<=(others=>'0');MULT_29<=((others=> (others=>'0')));
    SUM_PIXELS_30<=(others=>'0');MULT_30<=((others=> (others=>'0')));
    SUM_PIXELS_31<=(others=>'0');MULT_31<=((others=> (others=>'0')));
    SUM_PIXELS_32<=(others=>'0');MULT_32<=((others=> (others=>'0')));
    SUM_PIXELS_33<=(others=>'0');MULT_33<=((others=> (others=>'0')));
    SUM_PIXELS_34<=(others=>'0');MULT_34<=((others=> (others=>'0')));
    SUM_PIXELS_35<=(others=>'0');MULT_35<=((others=> (others=>'0')));
    SUM_PIXELS_36<=(others=>'0');MULT_36<=((others=> (others=>'0')));
    SUM_PIXELS_37<=(others=>'0');MULT_37<=((others=> (others=>'0')));
    SUM_PIXELS_38<=(others=>'0');MULT_38<=((others=> (others=>'0')));
    SUM_PIXELS_39<=(others=>'0');MULT_39<=((others=> (others=>'0')));
    SUM_PIXELS_40<=(others=>'0');MULT_40<=((others=> (others=>'0')));
    SUM_PIXELS_41<=(others=>'0');MULT_41<=((others=> (others=>'0')));
    SUM_PIXELS_42<=(others=>'0');MULT_42<=((others=> (others=>'0')));
    SUM_PIXELS_43<=(others=>'0');MULT_43<=((others=> (others=>'0')));
    SUM_PIXELS_44<=(others=>'0');MULT_44<=((others=> (others=>'0')));
    SUM_PIXELS_45<=(others=>'0');MULT_45<=((others=> (others=>'0')));
    SUM_PIXELS_46<=(others=>'0');MULT_46<=((others=> (others=>'0')));
    SUM_PIXELS_47<=(others=>'0');MULT_47<=((others=> (others=>'0')));
    SUM_PIXELS_48<=(others=>'0');MULT_48<=((others=> (others=>'0')));
    SUM_PIXELS_49<=(others=>'0');MULT_49<=((others=> (others=>'0')));
    SUM_PIXELS_50<=(others=>'0');MULT_50<=((others=> (others=>'0')));
    SUM_PIXELS_51<=(others=>'0');MULT_51<=((others=> (others=>'0')));
    SUM_PIXELS_52<=(others=>'0');MULT_52<=((others=> (others=>'0')));
    SUM_PIXELS_53<=(others=>'0');MULT_53<=((others=> (others=>'0')));
    SUM_PIXELS_54<=(others=>'0');MULT_54<=((others=> (others=>'0')));
    SUM_PIXELS_55<=(others=>'0');MULT_55<=((others=> (others=>'0')));
    SUM_PIXELS_56<=(others=>'0');MULT_56<=((others=> (others=>'0')));
    SUM_PIXELS_57<=(others=>'0');MULT_57<=((others=> (others=>'0')));
    SUM_PIXELS_58<=(others=>'0');MULT_58<=((others=> (others=>'0')));
    SUM_PIXELS_59<=(others=>'0');MULT_59<=((others=> (others=>'0')));
    SUM_PIXELS_60<=(others=>'0');MULT_60<=((others=> (others=>'0')));
    SUM_PIXELS_61<=(others=>'0');MULT_61<=((others=> (others=>'0')));
    SUM_PIXELS_62<=(others=>'0');MULT_62<=((others=> (others=>'0')));
    SUM_PIXELS_63<=(others=>'0');MULT_63<=((others=> (others=>'0')));
    SUM_PIXELS_64<=(others=>'0');MULT_64<=((others=> (others=>'0')));
    SUM_PIXELS_65<=(others=>'0');MULT_65<=((others=> (others=>'0')));
    SUM_PIXELS_66<=(others=>'0');MULT_66<=((others=> (others=>'0')));
    SUM_PIXELS_67<=(others=>'0');MULT_67<=((others=> (others=>'0')));
    SUM_PIXELS_68<=(others=>'0');MULT_68<=((others=> (others=>'0')));
    SUM_PIXELS_69<=(others=>'0');MULT_69<=((others=> (others=>'0')));
    SUM_PIXELS_70<=(others=>'0');MULT_70<=((others=> (others=>'0')));
    SUM_PIXELS_71<=(others=>'0');MULT_71<=((others=> (others=>'0')));
    SUM_PIXELS_72<=(others=>'0');MULT_72<=((others=> (others=>'0')));
    SUM_PIXELS_73<=(others=>'0');MULT_73<=((others=> (others=>'0')));
    SUM_PIXELS_74<=(others=>'0');MULT_74<=((others=> (others=>'0')));
    SUM_PIXELS_75<=(others=>'0');MULT_75<=((others=> (others=>'0')));
    SUM_PIXELS_76<=(others=>'0');MULT_76<=((others=> (others=>'0')));
    SUM_PIXELS_77<=(others=>'0');MULT_77<=((others=> (others=>'0')));
    SUM_PIXELS_78<=(others=>'0');MULT_78<=((others=> (others=>'0')));
    SUM_PIXELS_79<=(others=>'0');MULT_79<=((others=> (others=>'0')));
    SUM_PIXELS_80<=(others=>'0');MULT_80<=((others=> (others=>'0')));
    SUM_PIXELS_81<=(others=>'0');MULT_81<=((others=> (others=>'0')));
    SUM_PIXELS_82<=(others=>'0');MULT_82<=((others=> (others=>'0')));
    SUM_PIXELS_83<=(others=>'0');MULT_83<=((others=> (others=>'0')));
    SUM_PIXELS_84<=(others=>'0');MULT_84<=((others=> (others=>'0')));
    SUM_PIXELS_85<=(others=>'0');MULT_85<=((others=> (others=>'0')));
    SUM_PIXELS_86<=(others=>'0');MULT_86<=((others=> (others=>'0')));
    SUM_PIXELS_87<=(others=>'0');MULT_87<=((others=> (others=>'0')));
    SUM_PIXELS_88<=(others=>'0');MULT_88<=((others=> (others=>'0')));
    SUM_PIXELS_89<=(others=>'0');MULT_89<=((others=> (others=>'0')));
    SUM_PIXELS_90<=(others=>'0');MULT_90<=((others=> (others=>'0')));
    SUM_PIXELS_91<=(others=>'0');MULT_91<=((others=> (others=>'0')));
    SUM_PIXELS_92<=(others=>'0');MULT_92<=((others=> (others=>'0')));
    SUM_PIXELS_93<=(others=>'0');MULT_93<=((others=> (others=>'0')));
    SUM_PIXELS_94<=(others=>'0');MULT_94<=((others=> (others=>'0')));
    SUM_PIXELS_95<=(others=>'0');MULT_95<=((others=> (others=>'0')));
    SUM_PIXELS_96<=(others=>'0');MULT_96<=((others=> (others=>'0')));
    SUM_PIXELS_97<=(others=>'0');MULT_97<=((others=> (others=>'0')));
    SUM_PIXELS_98<=(others=>'0');MULT_98<=((others=> (others=>'0')));
    SUM_PIXELS_99<=(others=>'0');MULT_99<=((others=> (others=>'0')));
    SUM_PIXELS_100<=(others=>'0');MULT_100<=((others=> (others=>'0')));
    SUM_PIXELS_101<=(others=>'0');MULT_101<=((others=> (others=>'0')));
    SUM_PIXELS_102<=(others=>'0');MULT_102<=((others=> (others=>'0')));
    SUM_PIXELS_103<=(others=>'0');MULT_103<=((others=> (others=>'0')));
    SUM_PIXELS_104<=(others=>'0');MULT_104<=((others=> (others=>'0')));
    SUM_PIXELS_105<=(others=>'0');MULT_105<=((others=> (others=>'0')));
    SUM_PIXELS_106<=(others=>'0');MULT_106<=((others=> (others=>'0')));
    SUM_PIXELS_107<=(others=>'0');MULT_107<=((others=> (others=>'0')));
    SUM_PIXELS_108<=(others=>'0');MULT_108<=((others=> (others=>'0')));
    SUM_PIXELS_109<=(others=>'0');MULT_109<=((others=> (others=>'0')));
    SUM_PIXELS_110<=(others=>'0');MULT_110<=((others=> (others=>'0')));
    SUM_PIXELS_111<=(others=>'0');MULT_111<=((others=> (others=>'0')));
    SUM_PIXELS_112<=(others=>'0');MULT_112<=((others=> (others=>'0')));
    SUM_PIXELS_113<=(others=>'0');MULT_113<=((others=> (others=>'0')));
    SUM_PIXELS_114<=(others=>'0');MULT_114<=((others=> (others=>'0')));
    SUM_PIXELS_115<=(others=>'0');MULT_115<=((others=> (others=>'0')));
    SUM_PIXELS_116<=(others=>'0');MULT_116<=((others=> (others=>'0')));
    SUM_PIXELS_117<=(others=>'0');MULT_117<=((others=> (others=>'0')));
    SUM_PIXELS_118<=(others=>'0');MULT_118<=((others=> (others=>'0')));
    SUM_PIXELS_119<=(others=>'0');MULT_119<=((others=> (others=>'0')));
    SUM_PIXELS_120<=(others=>'0');MULT_120<=((others=> (others=>'0')));

    EN_SUM_MULT_1<='0';
    MULTS_1_1<=((others=> (others=>'0')));
    MULTS_1_2<=((others=> (others=>'0')));
    MULTS_1_3<=((others=> (others=>'0')));
    MULTS_1_4<=((others=> (others=>'0')));
    MULTS_1_5<=((others=> (others=>'0')));
    MULTS_1_6<=((others=> (others=>'0')));
    MULTS_1_7<=((others=> (others=>'0')));
    MULTS_1_8<=((others=> (others=>'0')));
    MULTS_1_9<=((others=> (others=>'0')));
    MULTS_1_10<=((others=> (others=>'0')));
    MULTS_1_11<=((others=> (others=>'0')));
    MULTS_1_12<=((others=> (others=>'0')));
    MULTS_1_13<=((others=> (others=>'0')));
    MULTS_1_14<=((others=> (others=>'0')));
    MULTS_1_15<=((others=> (others=>'0')));
    MULTS_1_16<=((others=> (others=>'0')));
    MULTS_1_17<=((others=> (others=>'0')));
    MULTS_1_18<=((others=> (others=>'0')));
    MULTS_1_19<=((others=> (others=>'0')));
    MULTS_1_20<=((others=> (others=>'0')));
    MULTS_1_21<=((others=> (others=>'0')));
    MULTS_1_22<=((others=> (others=>'0')));
    MULTS_1_23<=((others=> (others=>'0')));
    MULTS_1_24<=((others=> (others=>'0')));
    MULTS_1_25<=((others=> (others=>'0')));
    MULTS_1_26<=((others=> (others=>'0')));
    MULTS_1_27<=((others=> (others=>'0')));
    MULTS_1_28<=((others=> (others=>'0')));
    MULTS_1_29<=((others=> (others=>'0')));
    MULTS_1_30<=((others=> (others=>'0')));
    MULTS_1_31<=((others=> (others=>'0')));
    MULTS_1_32<=((others=> (others=>'0')));
    MULTS_1_33<=((others=> (others=>'0')));
    MULTS_1_34<=((others=> (others=>'0')));
    MULTS_1_35<=((others=> (others=>'0')));
    MULTS_1_36<=((others=> (others=>'0')));
    MULTS_1_37<=((others=> (others=>'0')));
    MULTS_1_38<=((others=> (others=>'0')));
    MULTS_1_39<=((others=> (others=>'0')));
    MULTS_1_40<=((others=> (others=>'0')));
    MULTS_1_41<=((others=> (others=>'0')));
    MULTS_1_42<=((others=> (others=>'0')));
    MULTS_1_43<=((others=> (others=>'0')));
    MULTS_1_44<=((others=> (others=>'0')));
    MULTS_1_45<=((others=> (others=>'0')));
    MULTS_1_46<=((others=> (others=>'0')));
    MULTS_1_47<=((others=> (others=>'0')));
    MULTS_1_48<=((others=> (others=>'0')));
    MULTS_1_49<=((others=> (others=>'0')));
    MULTS_1_50<=((others=> (others=>'0')));
    MULTS_1_51<=((others=> (others=>'0')));
    MULTS_1_52<=((others=> (others=>'0')));
    MULTS_1_53<=((others=> (others=>'0')));
    MULTS_1_54<=((others=> (others=>'0')));
    MULTS_1_55<=((others=> (others=>'0')));
    MULTS_1_56<=((others=> (others=>'0')));
    MULTS_1_57<=((others=> (others=>'0')));
    MULTS_1_58<=((others=> (others=>'0')));
    MULTS_1_59<=((others=> (others=>'0')));
    MULTS_1_60<=((others=> (others=>'0')));
    MULTS_1_61<=((others=> (others=>'0')));
    MULTS_1_62<=((others=> (others=>'0')));
    MULTS_1_63<=((others=> (others=>'0')));
    MULTS_1_64<=((others=> (others=>'0')));
    MULTS_1_65<=((others=> (others=>'0')));
    MULTS_1_66<=((others=> (others=>'0')));
    MULTS_1_67<=((others=> (others=>'0')));
    MULTS_1_68<=((others=> (others=>'0')));
    MULTS_1_69<=((others=> (others=>'0')));
    MULTS_1_70<=((others=> (others=>'0')));
    MULTS_1_71<=((others=> (others=>'0')));
    MULTS_1_72<=((others=> (others=>'0')));
    MULTS_1_73<=((others=> (others=>'0')));
    MULTS_1_74<=((others=> (others=>'0')));
    MULTS_1_75<=((others=> (others=>'0')));
    MULTS_1_76<=((others=> (others=>'0')));
    MULTS_1_77<=((others=> (others=>'0')));
    MULTS_1_78<=((others=> (others=>'0')));
    MULTS_1_79<=((others=> (others=>'0')));
    MULTS_1_80<=((others=> (others=>'0')));
    MULTS_1_81<=((others=> (others=>'0')));
    MULTS_1_82<=((others=> (others=>'0')));
    MULTS_1_83<=((others=> (others=>'0')));
    MULTS_1_84<=((others=> (others=>'0')));
    MULTS_1_85<=((others=> (others=>'0')));
    MULTS_1_86<=((others=> (others=>'0')));
    MULTS_1_87<=((others=> (others=>'0')));
    MULTS_1_88<=((others=> (others=>'0')));
    MULTS_1_89<=((others=> (others=>'0')));
    MULTS_1_90<=((others=> (others=>'0')));
    MULTS_1_91<=((others=> (others=>'0')));
    MULTS_1_92<=((others=> (others=>'0')));
    MULTS_1_93<=((others=> (others=>'0')));
    MULTS_1_94<=((others=> (others=>'0')));
    MULTS_1_95<=((others=> (others=>'0')));
    MULTS_1_96<=((others=> (others=>'0')));
    MULTS_1_97<=((others=> (others=>'0')));
    MULTS_1_98<=((others=> (others=>'0')));
    MULTS_1_99<=((others=> (others=>'0')));
    MULTS_1_100<=((others=> (others=>'0')));
    MULTS_1_101<=((others=> (others=>'0')));
    MULTS_1_102<=((others=> (others=>'0')));
    MULTS_1_103<=((others=> (others=>'0')));
    MULTS_1_104<=((others=> (others=>'0')));
    MULTS_1_105<=((others=> (others=>'0')));
    MULTS_1_106<=((others=> (others=>'0')));
    MULTS_1_107<=((others=> (others=>'0')));
    MULTS_1_108<=((others=> (others=>'0')));
    MULTS_1_109<=((others=> (others=>'0')));
    MULTS_1_110<=((others=> (others=>'0')));
    MULTS_1_111<=((others=> (others=>'0')));
    MULTS_1_112<=((others=> (others=>'0')));
    MULTS_1_113<=((others=> (others=>'0')));
    MULTS_1_114<=((others=> (others=>'0')));
    MULTS_1_115<=((others=> (others=>'0')));
    MULTS_1_116<=((others=> (others=>'0')));
    MULTS_1_117<=((others=> (others=>'0')));
    MULTS_1_118<=((others=> (others=>'0')));
    MULTS_1_119<=((others=> (others=>'0')));
    MULTS_1_120<=((others=> (others=>'0')));
    EN_SUM_MULT_2<='0';
    MULTS_2_1<=((others=> (others=>'0')));
    MULTS_2_2<=((others=> (others=>'0')));
    MULTS_2_3<=((others=> (others=>'0')));
    MULTS_2_4<=((others=> (others=>'0')));
    MULTS_2_5<=((others=> (others=>'0')));
    MULTS_2_6<=((others=> (others=>'0')));
    MULTS_2_7<=((others=> (others=>'0')));
    MULTS_2_8<=((others=> (others=>'0')));
    MULTS_2_9<=((others=> (others=>'0')));
    MULTS_2_10<=((others=> (others=>'0')));
    MULTS_2_11<=((others=> (others=>'0')));
    MULTS_2_12<=((others=> (others=>'0')));
    MULTS_2_13<=((others=> (others=>'0')));
    MULTS_2_14<=((others=> (others=>'0')));
    MULTS_2_15<=((others=> (others=>'0')));
    MULTS_2_16<=((others=> (others=>'0')));
    MULTS_2_17<=((others=> (others=>'0')));
    MULTS_2_18<=((others=> (others=>'0')));
    MULTS_2_19<=((others=> (others=>'0')));
    MULTS_2_20<=((others=> (others=>'0')));
    MULTS_2_21<=((others=> (others=>'0')));
    MULTS_2_22<=((others=> (others=>'0')));
    MULTS_2_23<=((others=> (others=>'0')));
    MULTS_2_24<=((others=> (others=>'0')));
    MULTS_2_25<=((others=> (others=>'0')));
    MULTS_2_26<=((others=> (others=>'0')));
    MULTS_2_27<=((others=> (others=>'0')));
    MULTS_2_28<=((others=> (others=>'0')));
    MULTS_2_29<=((others=> (others=>'0')));
    MULTS_2_30<=((others=> (others=>'0')));
    MULTS_2_31<=((others=> (others=>'0')));
    MULTS_2_32<=((others=> (others=>'0')));
    MULTS_2_33<=((others=> (others=>'0')));
    MULTS_2_34<=((others=> (others=>'0')));
    MULTS_2_35<=((others=> (others=>'0')));
    MULTS_2_36<=((others=> (others=>'0')));
    MULTS_2_37<=((others=> (others=>'0')));
    MULTS_2_38<=((others=> (others=>'0')));
    MULTS_2_39<=((others=> (others=>'0')));
    MULTS_2_40<=((others=> (others=>'0')));
    MULTS_2_41<=((others=> (others=>'0')));
    MULTS_2_42<=((others=> (others=>'0')));
    MULTS_2_43<=((others=> (others=>'0')));
    MULTS_2_44<=((others=> (others=>'0')));
    MULTS_2_45<=((others=> (others=>'0')));
    MULTS_2_46<=((others=> (others=>'0')));
    MULTS_2_47<=((others=> (others=>'0')));
    MULTS_2_48<=((others=> (others=>'0')));
    MULTS_2_49<=((others=> (others=>'0')));
    MULTS_2_50<=((others=> (others=>'0')));
    MULTS_2_51<=((others=> (others=>'0')));
    MULTS_2_52<=((others=> (others=>'0')));
    MULTS_2_53<=((others=> (others=>'0')));
    MULTS_2_54<=((others=> (others=>'0')));
    MULTS_2_55<=((others=> (others=>'0')));
    MULTS_2_56<=((others=> (others=>'0')));
    MULTS_2_57<=((others=> (others=>'0')));
    MULTS_2_58<=((others=> (others=>'0')));
    MULTS_2_59<=((others=> (others=>'0')));
    MULTS_2_60<=((others=> (others=>'0')));
    MULTS_2_61<=((others=> (others=>'0')));
    MULTS_2_62<=((others=> (others=>'0')));
    MULTS_2_63<=((others=> (others=>'0')));
    MULTS_2_64<=((others=> (others=>'0')));
    MULTS_2_65<=((others=> (others=>'0')));
    MULTS_2_66<=((others=> (others=>'0')));
    MULTS_2_67<=((others=> (others=>'0')));
    MULTS_2_68<=((others=> (others=>'0')));
    MULTS_2_69<=((others=> (others=>'0')));
    MULTS_2_70<=((others=> (others=>'0')));
    MULTS_2_71<=((others=> (others=>'0')));
    MULTS_2_72<=((others=> (others=>'0')));
    MULTS_2_73<=((others=> (others=>'0')));
    MULTS_2_74<=((others=> (others=>'0')));
    MULTS_2_75<=((others=> (others=>'0')));
    MULTS_2_76<=((others=> (others=>'0')));
    MULTS_2_77<=((others=> (others=>'0')));
    MULTS_2_78<=((others=> (others=>'0')));
    MULTS_2_79<=((others=> (others=>'0')));
    MULTS_2_80<=((others=> (others=>'0')));
    MULTS_2_81<=((others=> (others=>'0')));
    MULTS_2_82<=((others=> (others=>'0')));
    MULTS_2_83<=((others=> (others=>'0')));
    MULTS_2_84<=((others=> (others=>'0')));
    MULTS_2_85<=((others=> (others=>'0')));
    MULTS_2_86<=((others=> (others=>'0')));
    MULTS_2_87<=((others=> (others=>'0')));
    MULTS_2_88<=((others=> (others=>'0')));
    MULTS_2_89<=((others=> (others=>'0')));
    MULTS_2_90<=((others=> (others=>'0')));
    MULTS_2_91<=((others=> (others=>'0')));
    MULTS_2_92<=((others=> (others=>'0')));
    MULTS_2_93<=((others=> (others=>'0')));
    MULTS_2_94<=((others=> (others=>'0')));
    MULTS_2_95<=((others=> (others=>'0')));
    MULTS_2_96<=((others=> (others=>'0')));
    MULTS_2_97<=((others=> (others=>'0')));
    MULTS_2_98<=((others=> (others=>'0')));
    MULTS_2_99<=((others=> (others=>'0')));
    MULTS_2_100<=((others=> (others=>'0')));
    MULTS_2_101<=((others=> (others=>'0')));
    MULTS_2_102<=((others=> (others=>'0')));
    MULTS_2_103<=((others=> (others=>'0')));
    MULTS_2_104<=((others=> (others=>'0')));
    MULTS_2_105<=((others=> (others=>'0')));
    MULTS_2_106<=((others=> (others=>'0')));
    MULTS_2_107<=((others=> (others=>'0')));
    MULTS_2_108<=((others=> (others=>'0')));
    MULTS_2_109<=((others=> (others=>'0')));
    MULTS_2_110<=((others=> (others=>'0')));
    MULTS_2_111<=((others=> (others=>'0')));
    MULTS_2_112<=((others=> (others=>'0')));
    MULTS_2_113<=((others=> (others=>'0')));
    MULTS_2_114<=((others=> (others=>'0')));
    MULTS_2_115<=((others=> (others=>'0')));
    MULTS_2_116<=((others=> (others=>'0')));
    MULTS_2_117<=((others=> (others=>'0')));
    MULTS_2_118<=((others=> (others=>'0')));
    MULTS_2_119<=((others=> (others=>'0')));
    MULTS_2_120<=((others=> (others=>'0')));
    EN_SUM_MULT_3<='0';
    MULTS_3_1<=((others=> (others=>'0')));
    MULTS_3_2<=((others=> (others=>'0')));
    MULTS_3_3<=((others=> (others=>'0')));
    MULTS_3_4<=((others=> (others=>'0')));
    MULTS_3_5<=((others=> (others=>'0')));
    MULTS_3_6<=((others=> (others=>'0')));
    MULTS_3_7<=((others=> (others=>'0')));
    MULTS_3_8<=((others=> (others=>'0')));
    MULTS_3_9<=((others=> (others=>'0')));
    MULTS_3_10<=((others=> (others=>'0')));
    MULTS_3_11<=((others=> (others=>'0')));
    MULTS_3_12<=((others=> (others=>'0')));
    MULTS_3_13<=((others=> (others=>'0')));
    MULTS_3_14<=((others=> (others=>'0')));
    MULTS_3_15<=((others=> (others=>'0')));
    MULTS_3_16<=((others=> (others=>'0')));
    MULTS_3_17<=((others=> (others=>'0')));
    MULTS_3_18<=((others=> (others=>'0')));
    MULTS_3_19<=((others=> (others=>'0')));
    MULTS_3_20<=((others=> (others=>'0')));
    MULTS_3_21<=((others=> (others=>'0')));
    MULTS_3_22<=((others=> (others=>'0')));
    MULTS_3_23<=((others=> (others=>'0')));
    MULTS_3_24<=((others=> (others=>'0')));
    MULTS_3_25<=((others=> (others=>'0')));
    MULTS_3_26<=((others=> (others=>'0')));
    MULTS_3_27<=((others=> (others=>'0')));
    MULTS_3_28<=((others=> (others=>'0')));
    MULTS_3_29<=((others=> (others=>'0')));
    MULTS_3_30<=((others=> (others=>'0')));
    MULTS_3_31<=((others=> (others=>'0')));
    MULTS_3_32<=((others=> (others=>'0')));
    MULTS_3_33<=((others=> (others=>'0')));
    MULTS_3_34<=((others=> (others=>'0')));
    MULTS_3_35<=((others=> (others=>'0')));
    MULTS_3_36<=((others=> (others=>'0')));
    MULTS_3_37<=((others=> (others=>'0')));
    MULTS_3_38<=((others=> (others=>'0')));
    MULTS_3_39<=((others=> (others=>'0')));
    MULTS_3_40<=((others=> (others=>'0')));
    MULTS_3_41<=((others=> (others=>'0')));
    MULTS_3_42<=((others=> (others=>'0')));
    MULTS_3_43<=((others=> (others=>'0')));
    MULTS_3_44<=((others=> (others=>'0')));
    MULTS_3_45<=((others=> (others=>'0')));
    MULTS_3_46<=((others=> (others=>'0')));
    MULTS_3_47<=((others=> (others=>'0')));
    MULTS_3_48<=((others=> (others=>'0')));
    MULTS_3_49<=((others=> (others=>'0')));
    MULTS_3_50<=((others=> (others=>'0')));
    MULTS_3_51<=((others=> (others=>'0')));
    MULTS_3_52<=((others=> (others=>'0')));
    MULTS_3_53<=((others=> (others=>'0')));
    MULTS_3_54<=((others=> (others=>'0')));
    MULTS_3_55<=((others=> (others=>'0')));
    MULTS_3_56<=((others=> (others=>'0')));
    MULTS_3_57<=((others=> (others=>'0')));
    MULTS_3_58<=((others=> (others=>'0')));
    MULTS_3_59<=((others=> (others=>'0')));
    MULTS_3_60<=((others=> (others=>'0')));
    MULTS_3_61<=((others=> (others=>'0')));
    MULTS_3_62<=((others=> (others=>'0')));
    MULTS_3_63<=((others=> (others=>'0')));
    MULTS_3_64<=((others=> (others=>'0')));
    MULTS_3_65<=((others=> (others=>'0')));
    MULTS_3_66<=((others=> (others=>'0')));
    MULTS_3_67<=((others=> (others=>'0')));
    MULTS_3_68<=((others=> (others=>'0')));
    MULTS_3_69<=((others=> (others=>'0')));
    MULTS_3_70<=((others=> (others=>'0')));
    MULTS_3_71<=((others=> (others=>'0')));
    MULTS_3_72<=((others=> (others=>'0')));
    MULTS_3_73<=((others=> (others=>'0')));
    MULTS_3_74<=((others=> (others=>'0')));
    MULTS_3_75<=((others=> (others=>'0')));
    MULTS_3_76<=((others=> (others=>'0')));
    MULTS_3_77<=((others=> (others=>'0')));
    MULTS_3_78<=((others=> (others=>'0')));
    MULTS_3_79<=((others=> (others=>'0')));
    MULTS_3_80<=((others=> (others=>'0')));
    MULTS_3_81<=((others=> (others=>'0')));
    MULTS_3_82<=((others=> (others=>'0')));
    MULTS_3_83<=((others=> (others=>'0')));
    MULTS_3_84<=((others=> (others=>'0')));
    MULTS_3_85<=((others=> (others=>'0')));
    MULTS_3_86<=((others=> (others=>'0')));
    MULTS_3_87<=((others=> (others=>'0')));
    MULTS_3_88<=((others=> (others=>'0')));
    MULTS_3_89<=((others=> (others=>'0')));
    MULTS_3_90<=((others=> (others=>'0')));
    MULTS_3_91<=((others=> (others=>'0')));
    MULTS_3_92<=((others=> (others=>'0')));
    MULTS_3_93<=((others=> (others=>'0')));
    MULTS_3_94<=((others=> (others=>'0')));
    MULTS_3_95<=((others=> (others=>'0')));
    MULTS_3_96<=((others=> (others=>'0')));
    MULTS_3_97<=((others=> (others=>'0')));
    MULTS_3_98<=((others=> (others=>'0')));
    MULTS_3_99<=((others=> (others=>'0')));
    MULTS_3_100<=((others=> (others=>'0')));
    MULTS_3_101<=((others=> (others=>'0')));
    MULTS_3_102<=((others=> (others=>'0')));
    MULTS_3_103<=((others=> (others=>'0')));
    MULTS_3_104<=((others=> (others=>'0')));
    MULTS_3_105<=((others=> (others=>'0')));
    MULTS_3_106<=((others=> (others=>'0')));
    MULTS_3_107<=((others=> (others=>'0')));
    MULTS_3_108<=((others=> (others=>'0')));
    MULTS_3_109<=((others=> (others=>'0')));
    MULTS_3_110<=((others=> (others=>'0')));
    MULTS_3_111<=((others=> (others=>'0')));
    MULTS_3_112<=((others=> (others=>'0')));
    MULTS_3_113<=((others=> (others=>'0')));
    MULTS_3_114<=((others=> (others=>'0')));
    MULTS_3_115<=((others=> (others=>'0')));
    MULTS_3_116<=((others=> (others=>'0')));
    MULTS_3_117<=((others=> (others=>'0')));
    MULTS_3_118<=((others=> (others=>'0')));
    MULTS_3_119<=((others=> (others=>'0')));
    MULTS_3_120<=((others=> (others=>'0')));
    EN_SUM_MULT_4<='0';
    MULTS_4_1<=((others=> (others=>'0')));
    MULTS_4_2<=((others=> (others=>'0')));
    MULTS_4_3<=((others=> (others=>'0')));
    MULTS_4_4<=((others=> (others=>'0')));
    MULTS_4_5<=((others=> (others=>'0')));
    MULTS_4_6<=((others=> (others=>'0')));
    MULTS_4_7<=((others=> (others=>'0')));
    MULTS_4_8<=((others=> (others=>'0')));
    MULTS_4_9<=((others=> (others=>'0')));
    MULTS_4_10<=((others=> (others=>'0')));
    MULTS_4_11<=((others=> (others=>'0')));
    MULTS_4_12<=((others=> (others=>'0')));
    MULTS_4_13<=((others=> (others=>'0')));
    MULTS_4_14<=((others=> (others=>'0')));
    MULTS_4_15<=((others=> (others=>'0')));
    MULTS_4_16<=((others=> (others=>'0')));
    MULTS_4_17<=((others=> (others=>'0')));
    MULTS_4_18<=((others=> (others=>'0')));
    MULTS_4_19<=((others=> (others=>'0')));
    MULTS_4_20<=((others=> (others=>'0')));
    MULTS_4_21<=((others=> (others=>'0')));
    MULTS_4_22<=((others=> (others=>'0')));
    MULTS_4_23<=((others=> (others=>'0')));
    MULTS_4_24<=((others=> (others=>'0')));
    MULTS_4_25<=((others=> (others=>'0')));
    MULTS_4_26<=((others=> (others=>'0')));
    MULTS_4_27<=((others=> (others=>'0')));
    MULTS_4_28<=((others=> (others=>'0')));
    MULTS_4_29<=((others=> (others=>'0')));
    MULTS_4_30<=((others=> (others=>'0')));
    MULTS_4_31<=((others=> (others=>'0')));
    MULTS_4_32<=((others=> (others=>'0')));
    MULTS_4_33<=((others=> (others=>'0')));
    MULTS_4_34<=((others=> (others=>'0')));
    MULTS_4_35<=((others=> (others=>'0')));
    MULTS_4_36<=((others=> (others=>'0')));
    MULTS_4_37<=((others=> (others=>'0')));
    MULTS_4_38<=((others=> (others=>'0')));
    MULTS_4_39<=((others=> (others=>'0')));
    MULTS_4_40<=((others=> (others=>'0')));
    MULTS_4_41<=((others=> (others=>'0')));
    MULTS_4_42<=((others=> (others=>'0')));
    MULTS_4_43<=((others=> (others=>'0')));
    MULTS_4_44<=((others=> (others=>'0')));
    MULTS_4_45<=((others=> (others=>'0')));
    MULTS_4_46<=((others=> (others=>'0')));
    MULTS_4_47<=((others=> (others=>'0')));
    MULTS_4_48<=((others=> (others=>'0')));
    MULTS_4_49<=((others=> (others=>'0')));
    MULTS_4_50<=((others=> (others=>'0')));
    MULTS_4_51<=((others=> (others=>'0')));
    MULTS_4_52<=((others=> (others=>'0')));
    MULTS_4_53<=((others=> (others=>'0')));
    MULTS_4_54<=((others=> (others=>'0')));
    MULTS_4_55<=((others=> (others=>'0')));
    MULTS_4_56<=((others=> (others=>'0')));
    MULTS_4_57<=((others=> (others=>'0')));
    MULTS_4_58<=((others=> (others=>'0')));
    MULTS_4_59<=((others=> (others=>'0')));
    MULTS_4_60<=((others=> (others=>'0')));
    MULTS_4_61<=((others=> (others=>'0')));
    MULTS_4_62<=((others=> (others=>'0')));
    MULTS_4_63<=((others=> (others=>'0')));
    MULTS_4_64<=((others=> (others=>'0')));
    MULTS_4_65<=((others=> (others=>'0')));
    MULTS_4_66<=((others=> (others=>'0')));
    MULTS_4_67<=((others=> (others=>'0')));
    MULTS_4_68<=((others=> (others=>'0')));
    MULTS_4_69<=((others=> (others=>'0')));
    MULTS_4_70<=((others=> (others=>'0')));
    MULTS_4_71<=((others=> (others=>'0')));
    MULTS_4_72<=((others=> (others=>'0')));
    MULTS_4_73<=((others=> (others=>'0')));
    MULTS_4_74<=((others=> (others=>'0')));
    MULTS_4_75<=((others=> (others=>'0')));
    MULTS_4_76<=((others=> (others=>'0')));
    MULTS_4_77<=((others=> (others=>'0')));
    MULTS_4_78<=((others=> (others=>'0')));
    MULTS_4_79<=((others=> (others=>'0')));
    MULTS_4_80<=((others=> (others=>'0')));
    MULTS_4_81<=((others=> (others=>'0')));
    MULTS_4_82<=((others=> (others=>'0')));
    MULTS_4_83<=((others=> (others=>'0')));
    MULTS_4_84<=((others=> (others=>'0')));
    MULTS_4_85<=((others=> (others=>'0')));
    MULTS_4_86<=((others=> (others=>'0')));
    MULTS_4_87<=((others=> (others=>'0')));
    MULTS_4_88<=((others=> (others=>'0')));
    MULTS_4_89<=((others=> (others=>'0')));
    MULTS_4_90<=((others=> (others=>'0')));
    MULTS_4_91<=((others=> (others=>'0')));
    MULTS_4_92<=((others=> (others=>'0')));
    MULTS_4_93<=((others=> (others=>'0')));
    MULTS_4_94<=((others=> (others=>'0')));
    MULTS_4_95<=((others=> (others=>'0')));
    MULTS_4_96<=((others=> (others=>'0')));
    MULTS_4_97<=((others=> (others=>'0')));
    MULTS_4_98<=((others=> (others=>'0')));
    MULTS_4_99<=((others=> (others=>'0')));
    MULTS_4_100<=((others=> (others=>'0')));
    MULTS_4_101<=((others=> (others=>'0')));
    MULTS_4_102<=((others=> (others=>'0')));
    MULTS_4_103<=((others=> (others=>'0')));
    MULTS_4_104<=((others=> (others=>'0')));
    MULTS_4_105<=((others=> (others=>'0')));
    MULTS_4_106<=((others=> (others=>'0')));
    MULTS_4_107<=((others=> (others=>'0')));
    MULTS_4_108<=((others=> (others=>'0')));
    MULTS_4_109<=((others=> (others=>'0')));
    MULTS_4_110<=((others=> (others=>'0')));
    MULTS_4_111<=((others=> (others=>'0')));
    MULTS_4_112<=((others=> (others=>'0')));
    MULTS_4_113<=((others=> (others=>'0')));
    MULTS_4_114<=((others=> (others=>'0')));
    MULTS_4_115<=((others=> (others=>'0')));
    MULTS_4_116<=((others=> (others=>'0')));
    MULTS_4_117<=((others=> (others=>'0')));
    MULTS_4_118<=((others=> (others=>'0')));
    MULTS_4_119<=((others=> (others=>'0')));
    MULTS_4_120<=((others=> (others=>'0')));
    EN_SUM_MULT_5<='0';
    MULTS_5_1<=((others=> (others=>'0')));
    MULTS_5_2<=((others=> (others=>'0')));
    MULTS_5_3<=((others=> (others=>'0')));
    MULTS_5_4<=((others=> (others=>'0')));
    MULTS_5_5<=((others=> (others=>'0')));
    MULTS_5_6<=((others=> (others=>'0')));
    MULTS_5_7<=((others=> (others=>'0')));
    MULTS_5_8<=((others=> (others=>'0')));
    MULTS_5_9<=((others=> (others=>'0')));
    MULTS_5_10<=((others=> (others=>'0')));
    MULTS_5_11<=((others=> (others=>'0')));
    MULTS_5_12<=((others=> (others=>'0')));
    MULTS_5_13<=((others=> (others=>'0')));
    MULTS_5_14<=((others=> (others=>'0')));
    MULTS_5_15<=((others=> (others=>'0')));
    MULTS_5_16<=((others=> (others=>'0')));
    MULTS_5_17<=((others=> (others=>'0')));
    MULTS_5_18<=((others=> (others=>'0')));
    MULTS_5_19<=((others=> (others=>'0')));
    MULTS_5_20<=((others=> (others=>'0')));
    MULTS_5_21<=((others=> (others=>'0')));
    MULTS_5_22<=((others=> (others=>'0')));
    MULTS_5_23<=((others=> (others=>'0')));
    MULTS_5_24<=((others=> (others=>'0')));
    MULTS_5_25<=((others=> (others=>'0')));
    MULTS_5_26<=((others=> (others=>'0')));
    MULTS_5_27<=((others=> (others=>'0')));
    MULTS_5_28<=((others=> (others=>'0')));
    MULTS_5_29<=((others=> (others=>'0')));
    MULTS_5_30<=((others=> (others=>'0')));
    MULTS_5_31<=((others=> (others=>'0')));
    MULTS_5_32<=((others=> (others=>'0')));
    MULTS_5_33<=((others=> (others=>'0')));
    MULTS_5_34<=((others=> (others=>'0')));
    MULTS_5_35<=((others=> (others=>'0')));
    MULTS_5_36<=((others=> (others=>'0')));
    MULTS_5_37<=((others=> (others=>'0')));
    MULTS_5_38<=((others=> (others=>'0')));
    MULTS_5_39<=((others=> (others=>'0')));
    MULTS_5_40<=((others=> (others=>'0')));
    MULTS_5_41<=((others=> (others=>'0')));
    MULTS_5_42<=((others=> (others=>'0')));
    MULTS_5_43<=((others=> (others=>'0')));
    MULTS_5_44<=((others=> (others=>'0')));
    MULTS_5_45<=((others=> (others=>'0')));
    MULTS_5_46<=((others=> (others=>'0')));
    MULTS_5_47<=((others=> (others=>'0')));
    MULTS_5_48<=((others=> (others=>'0')));
    MULTS_5_49<=((others=> (others=>'0')));
    MULTS_5_50<=((others=> (others=>'0')));
    MULTS_5_51<=((others=> (others=>'0')));
    MULTS_5_52<=((others=> (others=>'0')));
    MULTS_5_53<=((others=> (others=>'0')));
    MULTS_5_54<=((others=> (others=>'0')));
    MULTS_5_55<=((others=> (others=>'0')));
    MULTS_5_56<=((others=> (others=>'0')));
    MULTS_5_57<=((others=> (others=>'0')));
    MULTS_5_58<=((others=> (others=>'0')));
    MULTS_5_59<=((others=> (others=>'0')));
    MULTS_5_60<=((others=> (others=>'0')));
    MULTS_5_61<=((others=> (others=>'0')));
    MULTS_5_62<=((others=> (others=>'0')));
    MULTS_5_63<=((others=> (others=>'0')));
    MULTS_5_64<=((others=> (others=>'0')));
    MULTS_5_65<=((others=> (others=>'0')));
    MULTS_5_66<=((others=> (others=>'0')));
    MULTS_5_67<=((others=> (others=>'0')));
    MULTS_5_68<=((others=> (others=>'0')));
    MULTS_5_69<=((others=> (others=>'0')));
    MULTS_5_70<=((others=> (others=>'0')));
    MULTS_5_71<=((others=> (others=>'0')));
    MULTS_5_72<=((others=> (others=>'0')));
    MULTS_5_73<=((others=> (others=>'0')));
    MULTS_5_74<=((others=> (others=>'0')));
    MULTS_5_75<=((others=> (others=>'0')));
    MULTS_5_76<=((others=> (others=>'0')));
    MULTS_5_77<=((others=> (others=>'0')));
    MULTS_5_78<=((others=> (others=>'0')));
    MULTS_5_79<=((others=> (others=>'0')));
    MULTS_5_80<=((others=> (others=>'0')));
    MULTS_5_81<=((others=> (others=>'0')));
    MULTS_5_82<=((others=> (others=>'0')));
    MULTS_5_83<=((others=> (others=>'0')));
    MULTS_5_84<=((others=> (others=>'0')));
    MULTS_5_85<=((others=> (others=>'0')));
    MULTS_5_86<=((others=> (others=>'0')));
    MULTS_5_87<=((others=> (others=>'0')));
    MULTS_5_88<=((others=> (others=>'0')));
    MULTS_5_89<=((others=> (others=>'0')));
    MULTS_5_90<=((others=> (others=>'0')));
    MULTS_5_91<=((others=> (others=>'0')));
    MULTS_5_92<=((others=> (others=>'0')));
    MULTS_5_93<=((others=> (others=>'0')));
    MULTS_5_94<=((others=> (others=>'0')));
    MULTS_5_95<=((others=> (others=>'0')));
    MULTS_5_96<=((others=> (others=>'0')));
    MULTS_5_97<=((others=> (others=>'0')));
    MULTS_5_98<=((others=> (others=>'0')));
    MULTS_5_99<=((others=> (others=>'0')));
    MULTS_5_100<=((others=> (others=>'0')));
    MULTS_5_101<=((others=> (others=>'0')));
    MULTS_5_102<=((others=> (others=>'0')));
    MULTS_5_103<=((others=> (others=>'0')));
    MULTS_5_104<=((others=> (others=>'0')));
    MULTS_5_105<=((others=> (others=>'0')));
    MULTS_5_106<=((others=> (others=>'0')));
    MULTS_5_107<=((others=> (others=>'0')));
    MULTS_5_108<=((others=> (others=>'0')));
    MULTS_5_109<=((others=> (others=>'0')));
    MULTS_5_110<=((others=> (others=>'0')));
    MULTS_5_111<=((others=> (others=>'0')));
    MULTS_5_112<=((others=> (others=>'0')));
    MULTS_5_113<=((others=> (others=>'0')));
    MULTS_5_114<=((others=> (others=>'0')));
    MULTS_5_115<=((others=> (others=>'0')));
    MULTS_5_116<=((others=> (others=>'0')));
    MULTS_5_117<=((others=> (others=>'0')));
    MULTS_5_118<=((others=> (others=>'0')));
    MULTS_5_119<=((others=> (others=>'0')));
    MULTS_5_120<=((others=> (others=>'0')));
    EN_SUM_MULT_6<='0';
    MULTS_6_1<=((others=> (others=>'0')));
    MULTS_6_2<=((others=> (others=>'0')));
    MULTS_6_3<=((others=> (others=>'0')));
    MULTS_6_4<=((others=> (others=>'0')));
    MULTS_6_5<=((others=> (others=>'0')));
    MULTS_6_6<=((others=> (others=>'0')));
    MULTS_6_7<=((others=> (others=>'0')));
    MULTS_6_8<=((others=> (others=>'0')));
    MULTS_6_9<=((others=> (others=>'0')));
    MULTS_6_10<=((others=> (others=>'0')));
    MULTS_6_11<=((others=> (others=>'0')));
    MULTS_6_12<=((others=> (others=>'0')));
    MULTS_6_13<=((others=> (others=>'0')));
    MULTS_6_14<=((others=> (others=>'0')));
    MULTS_6_15<=((others=> (others=>'0')));
    MULTS_6_16<=((others=> (others=>'0')));
    MULTS_6_17<=((others=> (others=>'0')));
    MULTS_6_18<=((others=> (others=>'0')));
    MULTS_6_19<=((others=> (others=>'0')));
    MULTS_6_20<=((others=> (others=>'0')));
    MULTS_6_21<=((others=> (others=>'0')));
    MULTS_6_22<=((others=> (others=>'0')));
    MULTS_6_23<=((others=> (others=>'0')));
    MULTS_6_24<=((others=> (others=>'0')));
    MULTS_6_25<=((others=> (others=>'0')));
    MULTS_6_26<=((others=> (others=>'0')));
    MULTS_6_27<=((others=> (others=>'0')));
    MULTS_6_28<=((others=> (others=>'0')));
    MULTS_6_29<=((others=> (others=>'0')));
    MULTS_6_30<=((others=> (others=>'0')));
    MULTS_6_31<=((others=> (others=>'0')));
    MULTS_6_32<=((others=> (others=>'0')));
    MULTS_6_33<=((others=> (others=>'0')));
    MULTS_6_34<=((others=> (others=>'0')));
    MULTS_6_35<=((others=> (others=>'0')));
    MULTS_6_36<=((others=> (others=>'0')));
    MULTS_6_37<=((others=> (others=>'0')));
    MULTS_6_38<=((others=> (others=>'0')));
    MULTS_6_39<=((others=> (others=>'0')));
    MULTS_6_40<=((others=> (others=>'0')));
    MULTS_6_41<=((others=> (others=>'0')));
    MULTS_6_42<=((others=> (others=>'0')));
    MULTS_6_43<=((others=> (others=>'0')));
    MULTS_6_44<=((others=> (others=>'0')));
    MULTS_6_45<=((others=> (others=>'0')));
    MULTS_6_46<=((others=> (others=>'0')));
    MULTS_6_47<=((others=> (others=>'0')));
    MULTS_6_48<=((others=> (others=>'0')));
    MULTS_6_49<=((others=> (others=>'0')));
    MULTS_6_50<=((others=> (others=>'0')));
    MULTS_6_51<=((others=> (others=>'0')));
    MULTS_6_52<=((others=> (others=>'0')));
    MULTS_6_53<=((others=> (others=>'0')));
    MULTS_6_54<=((others=> (others=>'0')));
    MULTS_6_55<=((others=> (others=>'0')));
    MULTS_6_56<=((others=> (others=>'0')));
    MULTS_6_57<=((others=> (others=>'0')));
    MULTS_6_58<=((others=> (others=>'0')));
    MULTS_6_59<=((others=> (others=>'0')));
    MULTS_6_60<=((others=> (others=>'0')));
    MULTS_6_61<=((others=> (others=>'0')));
    MULTS_6_62<=((others=> (others=>'0')));
    MULTS_6_63<=((others=> (others=>'0')));
    MULTS_6_64<=((others=> (others=>'0')));
    MULTS_6_65<=((others=> (others=>'0')));
    MULTS_6_66<=((others=> (others=>'0')));
    MULTS_6_67<=((others=> (others=>'0')));
    MULTS_6_68<=((others=> (others=>'0')));
    MULTS_6_69<=((others=> (others=>'0')));
    MULTS_6_70<=((others=> (others=>'0')));
    MULTS_6_71<=((others=> (others=>'0')));
    MULTS_6_72<=((others=> (others=>'0')));
    MULTS_6_73<=((others=> (others=>'0')));
    MULTS_6_74<=((others=> (others=>'0')));
    MULTS_6_75<=((others=> (others=>'0')));
    MULTS_6_76<=((others=> (others=>'0')));
    MULTS_6_77<=((others=> (others=>'0')));
    MULTS_6_78<=((others=> (others=>'0')));
    MULTS_6_79<=((others=> (others=>'0')));
    MULTS_6_80<=((others=> (others=>'0')));
    MULTS_6_81<=((others=> (others=>'0')));
    MULTS_6_82<=((others=> (others=>'0')));
    MULTS_6_83<=((others=> (others=>'0')));
    MULTS_6_84<=((others=> (others=>'0')));
    MULTS_6_85<=((others=> (others=>'0')));
    MULTS_6_86<=((others=> (others=>'0')));
    MULTS_6_87<=((others=> (others=>'0')));
    MULTS_6_88<=((others=> (others=>'0')));
    MULTS_6_89<=((others=> (others=>'0')));
    MULTS_6_90<=((others=> (others=>'0')));
    MULTS_6_91<=((others=> (others=>'0')));
    MULTS_6_92<=((others=> (others=>'0')));
    MULTS_6_93<=((others=> (others=>'0')));
    MULTS_6_94<=((others=> (others=>'0')));
    MULTS_6_95<=((others=> (others=>'0')));
    MULTS_6_96<=((others=> (others=>'0')));
    MULTS_6_97<=((others=> (others=>'0')));
    MULTS_6_98<=((others=> (others=>'0')));
    MULTS_6_99<=((others=> (others=>'0')));
    MULTS_6_100<=((others=> (others=>'0')));
    MULTS_6_101<=((others=> (others=>'0')));
    MULTS_6_102<=((others=> (others=>'0')));
    MULTS_6_103<=((others=> (others=>'0')));
    MULTS_6_104<=((others=> (others=>'0')));
    MULTS_6_105<=((others=> (others=>'0')));
    MULTS_6_106<=((others=> (others=>'0')));
    MULTS_6_107<=((others=> (others=>'0')));
    MULTS_6_108<=((others=> (others=>'0')));
    MULTS_6_109<=((others=> (others=>'0')));
    MULTS_6_110<=((others=> (others=>'0')));
    MULTS_6_111<=((others=> (others=>'0')));
    MULTS_6_112<=((others=> (others=>'0')));
    MULTS_6_113<=((others=> (others=>'0')));
    MULTS_6_114<=((others=> (others=>'0')));
    MULTS_6_115<=((others=> (others=>'0')));
    MULTS_6_116<=((others=> (others=>'0')));
    MULTS_6_117<=((others=> (others=>'0')));
    MULTS_6_118<=((others=> (others=>'0')));
    MULTS_6_119<=((others=> (others=>'0')));
    MULTS_6_120<=((others=> (others=>'0')));
    EN_SUM_MULT_7<='0';
    MULTS_7_1<=((others=> (others=>'0')));
    MULTS_7_2<=((others=> (others=>'0')));
    MULTS_7_3<=((others=> (others=>'0')));
    MULTS_7_4<=((others=> (others=>'0')));
    MULTS_7_5<=((others=> (others=>'0')));
    MULTS_7_6<=((others=> (others=>'0')));
    MULTS_7_7<=((others=> (others=>'0')));
    MULTS_7_8<=((others=> (others=>'0')));
    MULTS_7_9<=((others=> (others=>'0')));
    MULTS_7_10<=((others=> (others=>'0')));
    MULTS_7_11<=((others=> (others=>'0')));
    MULTS_7_12<=((others=> (others=>'0')));
    MULTS_7_13<=((others=> (others=>'0')));
    MULTS_7_14<=((others=> (others=>'0')));
    MULTS_7_15<=((others=> (others=>'0')));
    MULTS_7_16<=((others=> (others=>'0')));
    MULTS_7_17<=((others=> (others=>'0')));
    MULTS_7_18<=((others=> (others=>'0')));
    MULTS_7_19<=((others=> (others=>'0')));
    MULTS_7_20<=((others=> (others=>'0')));
    MULTS_7_21<=((others=> (others=>'0')));
    MULTS_7_22<=((others=> (others=>'0')));
    MULTS_7_23<=((others=> (others=>'0')));
    MULTS_7_24<=((others=> (others=>'0')));
    MULTS_7_25<=((others=> (others=>'0')));
    MULTS_7_26<=((others=> (others=>'0')));
    MULTS_7_27<=((others=> (others=>'0')));
    MULTS_7_28<=((others=> (others=>'0')));
    MULTS_7_29<=((others=> (others=>'0')));
    MULTS_7_30<=((others=> (others=>'0')));
    MULTS_7_31<=((others=> (others=>'0')));
    MULTS_7_32<=((others=> (others=>'0')));
    MULTS_7_33<=((others=> (others=>'0')));
    MULTS_7_34<=((others=> (others=>'0')));
    MULTS_7_35<=((others=> (others=>'0')));
    MULTS_7_36<=((others=> (others=>'0')));
    MULTS_7_37<=((others=> (others=>'0')));
    MULTS_7_38<=((others=> (others=>'0')));
    MULTS_7_39<=((others=> (others=>'0')));
    MULTS_7_40<=((others=> (others=>'0')));
    MULTS_7_41<=((others=> (others=>'0')));
    MULTS_7_42<=((others=> (others=>'0')));
    MULTS_7_43<=((others=> (others=>'0')));
    MULTS_7_44<=((others=> (others=>'0')));
    MULTS_7_45<=((others=> (others=>'0')));
    MULTS_7_46<=((others=> (others=>'0')));
    MULTS_7_47<=((others=> (others=>'0')));
    MULTS_7_48<=((others=> (others=>'0')));
    MULTS_7_49<=((others=> (others=>'0')));
    MULTS_7_50<=((others=> (others=>'0')));
    MULTS_7_51<=((others=> (others=>'0')));
    MULTS_7_52<=((others=> (others=>'0')));
    MULTS_7_53<=((others=> (others=>'0')));
    MULTS_7_54<=((others=> (others=>'0')));
    MULTS_7_55<=((others=> (others=>'0')));
    MULTS_7_56<=((others=> (others=>'0')));
    MULTS_7_57<=((others=> (others=>'0')));
    MULTS_7_58<=((others=> (others=>'0')));
    MULTS_7_59<=((others=> (others=>'0')));
    MULTS_7_60<=((others=> (others=>'0')));
    MULTS_7_61<=((others=> (others=>'0')));
    MULTS_7_62<=((others=> (others=>'0')));
    MULTS_7_63<=((others=> (others=>'0')));
    MULTS_7_64<=((others=> (others=>'0')));
    MULTS_7_65<=((others=> (others=>'0')));
    MULTS_7_66<=((others=> (others=>'0')));
    MULTS_7_67<=((others=> (others=>'0')));
    MULTS_7_68<=((others=> (others=>'0')));
    MULTS_7_69<=((others=> (others=>'0')));
    MULTS_7_70<=((others=> (others=>'0')));
    MULTS_7_71<=((others=> (others=>'0')));
    MULTS_7_72<=((others=> (others=>'0')));
    MULTS_7_73<=((others=> (others=>'0')));
    MULTS_7_74<=((others=> (others=>'0')));
    MULTS_7_75<=((others=> (others=>'0')));
    MULTS_7_76<=((others=> (others=>'0')));
    MULTS_7_77<=((others=> (others=>'0')));
    MULTS_7_78<=((others=> (others=>'0')));
    MULTS_7_79<=((others=> (others=>'0')));
    MULTS_7_80<=((others=> (others=>'0')));
    MULTS_7_81<=((others=> (others=>'0')));
    MULTS_7_82<=((others=> (others=>'0')));
    MULTS_7_83<=((others=> (others=>'0')));
    MULTS_7_84<=((others=> (others=>'0')));
    MULTS_7_85<=((others=> (others=>'0')));
    MULTS_7_86<=((others=> (others=>'0')));
    MULTS_7_87<=((others=> (others=>'0')));
    MULTS_7_88<=((others=> (others=>'0')));
    MULTS_7_89<=((others=> (others=>'0')));
    MULTS_7_90<=((others=> (others=>'0')));
    MULTS_7_91<=((others=> (others=>'0')));
    MULTS_7_92<=((others=> (others=>'0')));
    MULTS_7_93<=((others=> (others=>'0')));
    MULTS_7_94<=((others=> (others=>'0')));
    MULTS_7_95<=((others=> (others=>'0')));
    MULTS_7_96<=((others=> (others=>'0')));
    MULTS_7_97<=((others=> (others=>'0')));
    MULTS_7_98<=((others=> (others=>'0')));
    MULTS_7_99<=((others=> (others=>'0')));
    MULTS_7_100<=((others=> (others=>'0')));
    MULTS_7_101<=((others=> (others=>'0')));
    MULTS_7_102<=((others=> (others=>'0')));
    MULTS_7_103<=((others=> (others=>'0')));
    MULTS_7_104<=((others=> (others=>'0')));
    MULTS_7_105<=((others=> (others=>'0')));
    MULTS_7_106<=((others=> (others=>'0')));
    MULTS_7_107<=((others=> (others=>'0')));
    MULTS_7_108<=((others=> (others=>'0')));
    MULTS_7_109<=((others=> (others=>'0')));
    MULTS_7_110<=((others=> (others=>'0')));
    MULTS_7_111<=((others=> (others=>'0')));
    MULTS_7_112<=((others=> (others=>'0')));
    MULTS_7_113<=((others=> (others=>'0')));
    MULTS_7_114<=((others=> (others=>'0')));
    MULTS_7_115<=((others=> (others=>'0')));
    MULTS_7_116<=((others=> (others=>'0')));
    MULTS_7_117<=((others=> (others=>'0')));
    MULTS_7_118<=((others=> (others=>'0')));
    MULTS_7_119<=((others=> (others=>'0')));
    MULTS_7_120<=((others=> (others=>'0')));

------------------------------------------------ PROCESS START------------------------------------------------------
	  
   else 	
	if EN_LOC_STREAM_7='1' and EN_STREAM= '1' and OUT_PIXEL_COUNT<VALID_CYCLES  then    -- check valid data and enable stream
		
		if  FRST_TIM_EN_7='1' then EN_NXT_LYR_7<='1';end if;

			MULT_1(0)<=signed(DIN_1_7)*signed(FMAP_1_1);
			MULT_2(0)<=signed(DIN_2_7)*signed(FMAP_1_2);
			MULT_3(0)<=signed(DIN_3_7)*signed(FMAP_1_3);
			MULT_4(0)<=signed(DIN_4_7)*signed(FMAP_1_4);
			MULT_5(0)<=signed(DIN_5_7)*signed(FMAP_1_5);
			MULT_6(0)<=signed(DIN_6_7)*signed(FMAP_1_6);
			MULT_7(0)<=signed(DIN_7_7)*signed(FMAP_1_7);
			MULT_8(0)<=signed(DIN_8_7)*signed(FMAP_1_8);
			MULT_9(0)<=signed(DIN_9_7)*signed(FMAP_1_9);
			MULT_10(0)<=signed(DIN_10_7)*signed(FMAP_1_10);
			MULT_11(0)<=signed(DIN_11_7)*signed(FMAP_1_11);
			MULT_12(0)<=signed(DIN_12_7)*signed(FMAP_1_12);
			MULT_13(0)<=signed(DIN_13_7)*signed(FMAP_1_13);
			MULT_14(0)<=signed(DIN_14_7)*signed(FMAP_1_14);
			MULT_15(0)<=signed(DIN_15_7)*signed(FMAP_1_15);
			MULT_16(0)<=signed(DIN_16_7)*signed(FMAP_1_16);
			MULT_17(0)<=signed(DIN_17_7)*signed(FMAP_1_17);
			MULT_18(0)<=signed(DIN_18_7)*signed(FMAP_1_18);
			MULT_19(0)<=signed(DIN_19_7)*signed(FMAP_1_19);
			MULT_20(0)<=signed(DIN_20_7)*signed(FMAP_1_20);
			MULT_21(0)<=signed(DIN_21_7)*signed(FMAP_1_21);
			MULT_22(0)<=signed(DIN_22_7)*signed(FMAP_1_22);
			MULT_23(0)<=signed(DIN_23_7)*signed(FMAP_1_23);
			MULT_24(0)<=signed(DIN_24_7)*signed(FMAP_1_24);
			MULT_25(0)<=signed(DIN_25_7)*signed(FMAP_1_25);
			MULT_26(0)<=signed(DIN_26_7)*signed(FMAP_1_26);
			MULT_27(0)<=signed(DIN_27_7)*signed(FMAP_1_27);
			MULT_28(0)<=signed(DIN_28_7)*signed(FMAP_1_28);
			MULT_29(0)<=signed(DIN_29_7)*signed(FMAP_1_29);
			MULT_30(0)<=signed(DIN_30_7)*signed(FMAP_1_30);
			MULT_31(0)<=signed(DIN_31_7)*signed(FMAP_1_31);
			MULT_32(0)<=signed(DIN_32_7)*signed(FMAP_1_32);
			MULT_33(0)<=signed(DIN_33_7)*signed(FMAP_1_33);
			MULT_34(0)<=signed(DIN_34_7)*signed(FMAP_1_34);
			MULT_35(0)<=signed(DIN_35_7)*signed(FMAP_1_35);
			MULT_36(0)<=signed(DIN_36_7)*signed(FMAP_1_36);
			MULT_37(0)<=signed(DIN_37_7)*signed(FMAP_1_37);
			MULT_38(0)<=signed(DIN_38_7)*signed(FMAP_1_38);
			MULT_39(0)<=signed(DIN_39_7)*signed(FMAP_1_39);
			MULT_40(0)<=signed(DIN_40_7)*signed(FMAP_1_40);
			MULT_41(0)<=signed(DIN_41_7)*signed(FMAP_1_41);
			MULT_42(0)<=signed(DIN_42_7)*signed(FMAP_1_42);
			MULT_43(0)<=signed(DIN_43_7)*signed(FMAP_1_43);
			MULT_44(0)<=signed(DIN_44_7)*signed(FMAP_1_44);
			MULT_45(0)<=signed(DIN_45_7)*signed(FMAP_1_45);
			MULT_46(0)<=signed(DIN_46_7)*signed(FMAP_1_46);
			MULT_47(0)<=signed(DIN_47_7)*signed(FMAP_1_47);
			MULT_48(0)<=signed(DIN_48_7)*signed(FMAP_1_48);
			MULT_49(0)<=signed(DIN_49_7)*signed(FMAP_1_49);
			MULT_50(0)<=signed(DIN_50_7)*signed(FMAP_1_50);
			MULT_51(0)<=signed(DIN_51_7)*signed(FMAP_1_51);
			MULT_52(0)<=signed(DIN_52_7)*signed(FMAP_1_52);
			MULT_53(0)<=signed(DIN_53_7)*signed(FMAP_1_53);
			MULT_54(0)<=signed(DIN_54_7)*signed(FMAP_1_54);
			MULT_55(0)<=signed(DIN_55_7)*signed(FMAP_1_55);
			MULT_56(0)<=signed(DIN_56_7)*signed(FMAP_1_56);
			MULT_57(0)<=signed(DIN_57_7)*signed(FMAP_1_57);
			MULT_58(0)<=signed(DIN_58_7)*signed(FMAP_1_58);
			MULT_59(0)<=signed(DIN_59_7)*signed(FMAP_1_59);
			MULT_60(0)<=signed(DIN_60_7)*signed(FMAP_1_60);
			MULT_61(0)<=signed(DIN_61_7)*signed(FMAP_1_61);
			MULT_62(0)<=signed(DIN_62_7)*signed(FMAP_1_62);
			MULT_63(0)<=signed(DIN_63_7)*signed(FMAP_1_63);
			MULT_64(0)<=signed(DIN_64_7)*signed(FMAP_1_64);
			MULT_65(0)<=signed(DIN_65_7)*signed(FMAP_1_65);
			MULT_66(0)<=signed(DIN_66_7)*signed(FMAP_1_66);
			MULT_67(0)<=signed(DIN_67_7)*signed(FMAP_1_67);
			MULT_68(0)<=signed(DIN_68_7)*signed(FMAP_1_68);
			MULT_69(0)<=signed(DIN_69_7)*signed(FMAP_1_69);
			MULT_70(0)<=signed(DIN_70_7)*signed(FMAP_1_70);
			MULT_71(0)<=signed(DIN_71_7)*signed(FMAP_1_71);
			MULT_72(0)<=signed(DIN_72_7)*signed(FMAP_1_72);
			MULT_73(0)<=signed(DIN_73_7)*signed(FMAP_1_73);
			MULT_74(0)<=signed(DIN_74_7)*signed(FMAP_1_74);
			MULT_75(0)<=signed(DIN_75_7)*signed(FMAP_1_75);
			MULT_76(0)<=signed(DIN_76_7)*signed(FMAP_1_76);
			MULT_77(0)<=signed(DIN_77_7)*signed(FMAP_1_77);
			MULT_78(0)<=signed(DIN_78_7)*signed(FMAP_1_78);
			MULT_79(0)<=signed(DIN_79_7)*signed(FMAP_1_79);
			MULT_80(0)<=signed(DIN_80_7)*signed(FMAP_1_80);
			MULT_81(0)<=signed(DIN_81_7)*signed(FMAP_1_81);
			MULT_82(0)<=signed(DIN_82_7)*signed(FMAP_1_82);
			MULT_83(0)<=signed(DIN_83_7)*signed(FMAP_1_83);
			MULT_84(0)<=signed(DIN_84_7)*signed(FMAP_1_84);
			MULT_85(0)<=signed(DIN_85_7)*signed(FMAP_1_85);
			MULT_86(0)<=signed(DIN_86_7)*signed(FMAP_1_86);
			MULT_87(0)<=signed(DIN_87_7)*signed(FMAP_1_87);
			MULT_88(0)<=signed(DIN_88_7)*signed(FMAP_1_88);
			MULT_89(0)<=signed(DIN_89_7)*signed(FMAP_1_89);
			MULT_90(0)<=signed(DIN_90_7)*signed(FMAP_1_90);
			MULT_91(0)<=signed(DIN_91_7)*signed(FMAP_1_91);
			MULT_92(0)<=signed(DIN_92_7)*signed(FMAP_1_92);
			MULT_93(0)<=signed(DIN_93_7)*signed(FMAP_1_93);
			MULT_94(0)<=signed(DIN_94_7)*signed(FMAP_1_94);
			MULT_95(0)<=signed(DIN_95_7)*signed(FMAP_1_95);
			MULT_96(0)<=signed(DIN_96_7)*signed(FMAP_1_96);
			MULT_97(0)<=signed(DIN_97_7)*signed(FMAP_1_97);
			MULT_98(0)<=signed(DIN_98_7)*signed(FMAP_1_98);
			MULT_99(0)<=signed(DIN_99_7)*signed(FMAP_1_99);
			MULT_100(0)<=signed(DIN_100_7)*signed(FMAP_1_100);
			MULT_101(0)<=signed(DIN_101_7)*signed(FMAP_1_101);
			MULT_102(0)<=signed(DIN_102_7)*signed(FMAP_1_102);
			MULT_103(0)<=signed(DIN_103_7)*signed(FMAP_1_103);
			MULT_104(0)<=signed(DIN_104_7)*signed(FMAP_1_104);
			MULT_105(0)<=signed(DIN_105_7)*signed(FMAP_1_105);
			MULT_106(0)<=signed(DIN_106_7)*signed(FMAP_1_106);
			MULT_107(0)<=signed(DIN_107_7)*signed(FMAP_1_107);
			MULT_108(0)<=signed(DIN_108_7)*signed(FMAP_1_108);
			MULT_109(0)<=signed(DIN_109_7)*signed(FMAP_1_109);
			MULT_110(0)<=signed(DIN_110_7)*signed(FMAP_1_110);
			MULT_111(0)<=signed(DIN_111_7)*signed(FMAP_1_111);
			MULT_112(0)<=signed(DIN_112_7)*signed(FMAP_1_112);
			MULT_113(0)<=signed(DIN_113_7)*signed(FMAP_1_113);
			MULT_114(0)<=signed(DIN_114_7)*signed(FMAP_1_114);
			MULT_115(0)<=signed(DIN_115_7)*signed(FMAP_1_115);
			MULT_116(0)<=signed(DIN_116_7)*signed(FMAP_1_116);
			MULT_117(0)<=signed(DIN_117_7)*signed(FMAP_1_117);
			MULT_118(0)<=signed(DIN_118_7)*signed(FMAP_1_118);
			MULT_119(0)<=signed(DIN_119_7)*signed(FMAP_1_119);
			MULT_120(0)<=signed(DIN_120_7)*signed(FMAP_1_120);

			MULT_1(1)<=signed(DIN_1_7)*signed(FMAP_2_1);
			MULT_2(1)<=signed(DIN_2_7)*signed(FMAP_2_2);
			MULT_3(1)<=signed(DIN_3_7)*signed(FMAP_2_3);
			MULT_4(1)<=signed(DIN_4_7)*signed(FMAP_2_4);
			MULT_5(1)<=signed(DIN_5_7)*signed(FMAP_2_5);
			MULT_6(1)<=signed(DIN_6_7)*signed(FMAP_2_6);
			MULT_7(1)<=signed(DIN_7_7)*signed(FMAP_2_7);
			MULT_8(1)<=signed(DIN_8_7)*signed(FMAP_2_8);
			MULT_9(1)<=signed(DIN_9_7)*signed(FMAP_2_9);
			MULT_10(1)<=signed(DIN_10_7)*signed(FMAP_2_10);
			MULT_11(1)<=signed(DIN_11_7)*signed(FMAP_2_11);
			MULT_12(1)<=signed(DIN_12_7)*signed(FMAP_2_12);
			MULT_13(1)<=signed(DIN_13_7)*signed(FMAP_2_13);
			MULT_14(1)<=signed(DIN_14_7)*signed(FMAP_2_14);
			MULT_15(1)<=signed(DIN_15_7)*signed(FMAP_2_15);
			MULT_16(1)<=signed(DIN_16_7)*signed(FMAP_2_16);
			MULT_17(1)<=signed(DIN_17_7)*signed(FMAP_2_17);
			MULT_18(1)<=signed(DIN_18_7)*signed(FMAP_2_18);
			MULT_19(1)<=signed(DIN_19_7)*signed(FMAP_2_19);
			MULT_20(1)<=signed(DIN_20_7)*signed(FMAP_2_20);
			MULT_21(1)<=signed(DIN_21_7)*signed(FMAP_2_21);
			MULT_22(1)<=signed(DIN_22_7)*signed(FMAP_2_22);
			MULT_23(1)<=signed(DIN_23_7)*signed(FMAP_2_23);
			MULT_24(1)<=signed(DIN_24_7)*signed(FMAP_2_24);
			MULT_25(1)<=signed(DIN_25_7)*signed(FMAP_2_25);
			MULT_26(1)<=signed(DIN_26_7)*signed(FMAP_2_26);
			MULT_27(1)<=signed(DIN_27_7)*signed(FMAP_2_27);
			MULT_28(1)<=signed(DIN_28_7)*signed(FMAP_2_28);
			MULT_29(1)<=signed(DIN_29_7)*signed(FMAP_2_29);
			MULT_30(1)<=signed(DIN_30_7)*signed(FMAP_2_30);
			MULT_31(1)<=signed(DIN_31_7)*signed(FMAP_2_31);
			MULT_32(1)<=signed(DIN_32_7)*signed(FMAP_2_32);
			MULT_33(1)<=signed(DIN_33_7)*signed(FMAP_2_33);
			MULT_34(1)<=signed(DIN_34_7)*signed(FMAP_2_34);
			MULT_35(1)<=signed(DIN_35_7)*signed(FMAP_2_35);
			MULT_36(1)<=signed(DIN_36_7)*signed(FMAP_2_36);
			MULT_37(1)<=signed(DIN_37_7)*signed(FMAP_2_37);
			MULT_38(1)<=signed(DIN_38_7)*signed(FMAP_2_38);
			MULT_39(1)<=signed(DIN_39_7)*signed(FMAP_2_39);
			MULT_40(1)<=signed(DIN_40_7)*signed(FMAP_2_40);
			MULT_41(1)<=signed(DIN_41_7)*signed(FMAP_2_41);
			MULT_42(1)<=signed(DIN_42_7)*signed(FMAP_2_42);
			MULT_43(1)<=signed(DIN_43_7)*signed(FMAP_2_43);
			MULT_44(1)<=signed(DIN_44_7)*signed(FMAP_2_44);
			MULT_45(1)<=signed(DIN_45_7)*signed(FMAP_2_45);
			MULT_46(1)<=signed(DIN_46_7)*signed(FMAP_2_46);
			MULT_47(1)<=signed(DIN_47_7)*signed(FMAP_2_47);
			MULT_48(1)<=signed(DIN_48_7)*signed(FMAP_2_48);
			MULT_49(1)<=signed(DIN_49_7)*signed(FMAP_2_49);
			MULT_50(1)<=signed(DIN_50_7)*signed(FMAP_2_50);
			MULT_51(1)<=signed(DIN_51_7)*signed(FMAP_2_51);
			MULT_52(1)<=signed(DIN_52_7)*signed(FMAP_2_52);
			MULT_53(1)<=signed(DIN_53_7)*signed(FMAP_2_53);
			MULT_54(1)<=signed(DIN_54_7)*signed(FMAP_2_54);
			MULT_55(1)<=signed(DIN_55_7)*signed(FMAP_2_55);
			MULT_56(1)<=signed(DIN_56_7)*signed(FMAP_2_56);
			MULT_57(1)<=signed(DIN_57_7)*signed(FMAP_2_57);
			MULT_58(1)<=signed(DIN_58_7)*signed(FMAP_2_58);
			MULT_59(1)<=signed(DIN_59_7)*signed(FMAP_2_59);
			MULT_60(1)<=signed(DIN_60_7)*signed(FMAP_2_60);
			MULT_61(1)<=signed(DIN_61_7)*signed(FMAP_2_61);
			MULT_62(1)<=signed(DIN_62_7)*signed(FMAP_2_62);
			MULT_63(1)<=signed(DIN_63_7)*signed(FMAP_2_63);
			MULT_64(1)<=signed(DIN_64_7)*signed(FMAP_2_64);
			MULT_65(1)<=signed(DIN_65_7)*signed(FMAP_2_65);
			MULT_66(1)<=signed(DIN_66_7)*signed(FMAP_2_66);
			MULT_67(1)<=signed(DIN_67_7)*signed(FMAP_2_67);
			MULT_68(1)<=signed(DIN_68_7)*signed(FMAP_2_68);
			MULT_69(1)<=signed(DIN_69_7)*signed(FMAP_2_69);
			MULT_70(1)<=signed(DIN_70_7)*signed(FMAP_2_70);
			MULT_71(1)<=signed(DIN_71_7)*signed(FMAP_2_71);
			MULT_72(1)<=signed(DIN_72_7)*signed(FMAP_2_72);
			MULT_73(1)<=signed(DIN_73_7)*signed(FMAP_2_73);
			MULT_74(1)<=signed(DIN_74_7)*signed(FMAP_2_74);
			MULT_75(1)<=signed(DIN_75_7)*signed(FMAP_2_75);
			MULT_76(1)<=signed(DIN_76_7)*signed(FMAP_2_76);
			MULT_77(1)<=signed(DIN_77_7)*signed(FMAP_2_77);
			MULT_78(1)<=signed(DIN_78_7)*signed(FMAP_2_78);
			MULT_79(1)<=signed(DIN_79_7)*signed(FMAP_2_79);
			MULT_80(1)<=signed(DIN_80_7)*signed(FMAP_2_80);
			MULT_81(1)<=signed(DIN_81_7)*signed(FMAP_2_81);
			MULT_82(1)<=signed(DIN_82_7)*signed(FMAP_2_82);
			MULT_83(1)<=signed(DIN_83_7)*signed(FMAP_2_83);
			MULT_84(1)<=signed(DIN_84_7)*signed(FMAP_2_84);
			MULT_85(1)<=signed(DIN_85_7)*signed(FMAP_2_85);
			MULT_86(1)<=signed(DIN_86_7)*signed(FMAP_2_86);
			MULT_87(1)<=signed(DIN_87_7)*signed(FMAP_2_87);
			MULT_88(1)<=signed(DIN_88_7)*signed(FMAP_2_88);
			MULT_89(1)<=signed(DIN_89_7)*signed(FMAP_2_89);
			MULT_90(1)<=signed(DIN_90_7)*signed(FMAP_2_90);
			MULT_91(1)<=signed(DIN_91_7)*signed(FMAP_2_91);
			MULT_92(1)<=signed(DIN_92_7)*signed(FMAP_2_92);
			MULT_93(1)<=signed(DIN_93_7)*signed(FMAP_2_93);
			MULT_94(1)<=signed(DIN_94_7)*signed(FMAP_2_94);
			MULT_95(1)<=signed(DIN_95_7)*signed(FMAP_2_95);
			MULT_96(1)<=signed(DIN_96_7)*signed(FMAP_2_96);
			MULT_97(1)<=signed(DIN_97_7)*signed(FMAP_2_97);
			MULT_98(1)<=signed(DIN_98_7)*signed(FMAP_2_98);
			MULT_99(1)<=signed(DIN_99_7)*signed(FMAP_2_99);
			MULT_100(1)<=signed(DIN_100_7)*signed(FMAP_2_100);
			MULT_101(1)<=signed(DIN_101_7)*signed(FMAP_2_101);
			MULT_102(1)<=signed(DIN_102_7)*signed(FMAP_2_102);
			MULT_103(1)<=signed(DIN_103_7)*signed(FMAP_2_103);
			MULT_104(1)<=signed(DIN_104_7)*signed(FMAP_2_104);
			MULT_105(1)<=signed(DIN_105_7)*signed(FMAP_2_105);
			MULT_106(1)<=signed(DIN_106_7)*signed(FMAP_2_106);
			MULT_107(1)<=signed(DIN_107_7)*signed(FMAP_2_107);
			MULT_108(1)<=signed(DIN_108_7)*signed(FMAP_2_108);
			MULT_109(1)<=signed(DIN_109_7)*signed(FMAP_2_109);
			MULT_110(1)<=signed(DIN_110_7)*signed(FMAP_2_110);
			MULT_111(1)<=signed(DIN_111_7)*signed(FMAP_2_111);
			MULT_112(1)<=signed(DIN_112_7)*signed(FMAP_2_112);
			MULT_113(1)<=signed(DIN_113_7)*signed(FMAP_2_113);
			MULT_114(1)<=signed(DIN_114_7)*signed(FMAP_2_114);
			MULT_115(1)<=signed(DIN_115_7)*signed(FMAP_2_115);
			MULT_116(1)<=signed(DIN_116_7)*signed(FMAP_2_116);
			MULT_117(1)<=signed(DIN_117_7)*signed(FMAP_2_117);
			MULT_118(1)<=signed(DIN_118_7)*signed(FMAP_2_118);
			MULT_119(1)<=signed(DIN_119_7)*signed(FMAP_2_119);
			MULT_120(1)<=signed(DIN_120_7)*signed(FMAP_2_120);

			MULT_1(2)<=signed(DIN_1_7)*signed(FMAP_3_1);
			MULT_2(2)<=signed(DIN_2_7)*signed(FMAP_3_2);
			MULT_3(2)<=signed(DIN_3_7)*signed(FMAP_3_3);
			MULT_4(2)<=signed(DIN_4_7)*signed(FMAP_3_4);
			MULT_5(2)<=signed(DIN_5_7)*signed(FMAP_3_5);
			MULT_6(2)<=signed(DIN_6_7)*signed(FMAP_3_6);
			MULT_7(2)<=signed(DIN_7_7)*signed(FMAP_3_7);
			MULT_8(2)<=signed(DIN_8_7)*signed(FMAP_3_8);
			MULT_9(2)<=signed(DIN_9_7)*signed(FMAP_3_9);
			MULT_10(2)<=signed(DIN_10_7)*signed(FMAP_3_10);
			MULT_11(2)<=signed(DIN_11_7)*signed(FMAP_3_11);
			MULT_12(2)<=signed(DIN_12_7)*signed(FMAP_3_12);
			MULT_13(2)<=signed(DIN_13_7)*signed(FMAP_3_13);
			MULT_14(2)<=signed(DIN_14_7)*signed(FMAP_3_14);
			MULT_15(2)<=signed(DIN_15_7)*signed(FMAP_3_15);
			MULT_16(2)<=signed(DIN_16_7)*signed(FMAP_3_16);
			MULT_17(2)<=signed(DIN_17_7)*signed(FMAP_3_17);
			MULT_18(2)<=signed(DIN_18_7)*signed(FMAP_3_18);
			MULT_19(2)<=signed(DIN_19_7)*signed(FMAP_3_19);
			MULT_20(2)<=signed(DIN_20_7)*signed(FMAP_3_20);
			MULT_21(2)<=signed(DIN_21_7)*signed(FMAP_3_21);
			MULT_22(2)<=signed(DIN_22_7)*signed(FMAP_3_22);
			MULT_23(2)<=signed(DIN_23_7)*signed(FMAP_3_23);
			MULT_24(2)<=signed(DIN_24_7)*signed(FMAP_3_24);
			MULT_25(2)<=signed(DIN_25_7)*signed(FMAP_3_25);
			MULT_26(2)<=signed(DIN_26_7)*signed(FMAP_3_26);
			MULT_27(2)<=signed(DIN_27_7)*signed(FMAP_3_27);
			MULT_28(2)<=signed(DIN_28_7)*signed(FMAP_3_28);
			MULT_29(2)<=signed(DIN_29_7)*signed(FMAP_3_29);
			MULT_30(2)<=signed(DIN_30_7)*signed(FMAP_3_30);
			MULT_31(2)<=signed(DIN_31_7)*signed(FMAP_3_31);
			MULT_32(2)<=signed(DIN_32_7)*signed(FMAP_3_32);
			MULT_33(2)<=signed(DIN_33_7)*signed(FMAP_3_33);
			MULT_34(2)<=signed(DIN_34_7)*signed(FMAP_3_34);
			MULT_35(2)<=signed(DIN_35_7)*signed(FMAP_3_35);
			MULT_36(2)<=signed(DIN_36_7)*signed(FMAP_3_36);
			MULT_37(2)<=signed(DIN_37_7)*signed(FMAP_3_37);
			MULT_38(2)<=signed(DIN_38_7)*signed(FMAP_3_38);
			MULT_39(2)<=signed(DIN_39_7)*signed(FMAP_3_39);
			MULT_40(2)<=signed(DIN_40_7)*signed(FMAP_3_40);
			MULT_41(2)<=signed(DIN_41_7)*signed(FMAP_3_41);
			MULT_42(2)<=signed(DIN_42_7)*signed(FMAP_3_42);
			MULT_43(2)<=signed(DIN_43_7)*signed(FMAP_3_43);
			MULT_44(2)<=signed(DIN_44_7)*signed(FMAP_3_44);
			MULT_45(2)<=signed(DIN_45_7)*signed(FMAP_3_45);
			MULT_46(2)<=signed(DIN_46_7)*signed(FMAP_3_46);
			MULT_47(2)<=signed(DIN_47_7)*signed(FMAP_3_47);
			MULT_48(2)<=signed(DIN_48_7)*signed(FMAP_3_48);
			MULT_49(2)<=signed(DIN_49_7)*signed(FMAP_3_49);
			MULT_50(2)<=signed(DIN_50_7)*signed(FMAP_3_50);
			MULT_51(2)<=signed(DIN_51_7)*signed(FMAP_3_51);
			MULT_52(2)<=signed(DIN_52_7)*signed(FMAP_3_52);
			MULT_53(2)<=signed(DIN_53_7)*signed(FMAP_3_53);
			MULT_54(2)<=signed(DIN_54_7)*signed(FMAP_3_54);
			MULT_55(2)<=signed(DIN_55_7)*signed(FMAP_3_55);
			MULT_56(2)<=signed(DIN_56_7)*signed(FMAP_3_56);
			MULT_57(2)<=signed(DIN_57_7)*signed(FMAP_3_57);
			MULT_58(2)<=signed(DIN_58_7)*signed(FMAP_3_58);
			MULT_59(2)<=signed(DIN_59_7)*signed(FMAP_3_59);
			MULT_60(2)<=signed(DIN_60_7)*signed(FMAP_3_60);
			MULT_61(2)<=signed(DIN_61_7)*signed(FMAP_3_61);
			MULT_62(2)<=signed(DIN_62_7)*signed(FMAP_3_62);
			MULT_63(2)<=signed(DIN_63_7)*signed(FMAP_3_63);
			MULT_64(2)<=signed(DIN_64_7)*signed(FMAP_3_64);
			MULT_65(2)<=signed(DIN_65_7)*signed(FMAP_3_65);
			MULT_66(2)<=signed(DIN_66_7)*signed(FMAP_3_66);
			MULT_67(2)<=signed(DIN_67_7)*signed(FMAP_3_67);
			MULT_68(2)<=signed(DIN_68_7)*signed(FMAP_3_68);
			MULT_69(2)<=signed(DIN_69_7)*signed(FMAP_3_69);
			MULT_70(2)<=signed(DIN_70_7)*signed(FMAP_3_70);
			MULT_71(2)<=signed(DIN_71_7)*signed(FMAP_3_71);
			MULT_72(2)<=signed(DIN_72_7)*signed(FMAP_3_72);
			MULT_73(2)<=signed(DIN_73_7)*signed(FMAP_3_73);
			MULT_74(2)<=signed(DIN_74_7)*signed(FMAP_3_74);
			MULT_75(2)<=signed(DIN_75_7)*signed(FMAP_3_75);
			MULT_76(2)<=signed(DIN_76_7)*signed(FMAP_3_76);
			MULT_77(2)<=signed(DIN_77_7)*signed(FMAP_3_77);
			MULT_78(2)<=signed(DIN_78_7)*signed(FMAP_3_78);
			MULT_79(2)<=signed(DIN_79_7)*signed(FMAP_3_79);
			MULT_80(2)<=signed(DIN_80_7)*signed(FMAP_3_80);
			MULT_81(2)<=signed(DIN_81_7)*signed(FMAP_3_81);
			MULT_82(2)<=signed(DIN_82_7)*signed(FMAP_3_82);
			MULT_83(2)<=signed(DIN_83_7)*signed(FMAP_3_83);
			MULT_84(2)<=signed(DIN_84_7)*signed(FMAP_3_84);
			MULT_85(2)<=signed(DIN_85_7)*signed(FMAP_3_85);
			MULT_86(2)<=signed(DIN_86_7)*signed(FMAP_3_86);
			MULT_87(2)<=signed(DIN_87_7)*signed(FMAP_3_87);
			MULT_88(2)<=signed(DIN_88_7)*signed(FMAP_3_88);
			MULT_89(2)<=signed(DIN_89_7)*signed(FMAP_3_89);
			MULT_90(2)<=signed(DIN_90_7)*signed(FMAP_3_90);
			MULT_91(2)<=signed(DIN_91_7)*signed(FMAP_3_91);
			MULT_92(2)<=signed(DIN_92_7)*signed(FMAP_3_92);
			MULT_93(2)<=signed(DIN_93_7)*signed(FMAP_3_93);
			MULT_94(2)<=signed(DIN_94_7)*signed(FMAP_3_94);
			MULT_95(2)<=signed(DIN_95_7)*signed(FMAP_3_95);
			MULT_96(2)<=signed(DIN_96_7)*signed(FMAP_3_96);
			MULT_97(2)<=signed(DIN_97_7)*signed(FMAP_3_97);
			MULT_98(2)<=signed(DIN_98_7)*signed(FMAP_3_98);
			MULT_99(2)<=signed(DIN_99_7)*signed(FMAP_3_99);
			MULT_100(2)<=signed(DIN_100_7)*signed(FMAP_3_100);
			MULT_101(2)<=signed(DIN_101_7)*signed(FMAP_3_101);
			MULT_102(2)<=signed(DIN_102_7)*signed(FMAP_3_102);
			MULT_103(2)<=signed(DIN_103_7)*signed(FMAP_3_103);
			MULT_104(2)<=signed(DIN_104_7)*signed(FMAP_3_104);
			MULT_105(2)<=signed(DIN_105_7)*signed(FMAP_3_105);
			MULT_106(2)<=signed(DIN_106_7)*signed(FMAP_3_106);
			MULT_107(2)<=signed(DIN_107_7)*signed(FMAP_3_107);
			MULT_108(2)<=signed(DIN_108_7)*signed(FMAP_3_108);
			MULT_109(2)<=signed(DIN_109_7)*signed(FMAP_3_109);
			MULT_110(2)<=signed(DIN_110_7)*signed(FMAP_3_110);
			MULT_111(2)<=signed(DIN_111_7)*signed(FMAP_3_111);
			MULT_112(2)<=signed(DIN_112_7)*signed(FMAP_3_112);
			MULT_113(2)<=signed(DIN_113_7)*signed(FMAP_3_113);
			MULT_114(2)<=signed(DIN_114_7)*signed(FMAP_3_114);
			MULT_115(2)<=signed(DIN_115_7)*signed(FMAP_3_115);
			MULT_116(2)<=signed(DIN_116_7)*signed(FMAP_3_116);
			MULT_117(2)<=signed(DIN_117_7)*signed(FMAP_3_117);
			MULT_118(2)<=signed(DIN_118_7)*signed(FMAP_3_118);
			MULT_119(2)<=signed(DIN_119_7)*signed(FMAP_3_119);
			MULT_120(2)<=signed(DIN_120_7)*signed(FMAP_3_120);

			MULT_1(3)<=signed(DIN_1_7)*signed(FMAP_4_1);
			MULT_2(3)<=signed(DIN_2_7)*signed(FMAP_4_2);
			MULT_3(3)<=signed(DIN_3_7)*signed(FMAP_4_3);
			MULT_4(3)<=signed(DIN_4_7)*signed(FMAP_4_4);
			MULT_5(3)<=signed(DIN_5_7)*signed(FMAP_4_5);
			MULT_6(3)<=signed(DIN_6_7)*signed(FMAP_4_6);
			MULT_7(3)<=signed(DIN_7_7)*signed(FMAP_4_7);
			MULT_8(3)<=signed(DIN_8_7)*signed(FMAP_4_8);
			MULT_9(3)<=signed(DIN_9_7)*signed(FMAP_4_9);
			MULT_10(3)<=signed(DIN_10_7)*signed(FMAP_4_10);
			MULT_11(3)<=signed(DIN_11_7)*signed(FMAP_4_11);
			MULT_12(3)<=signed(DIN_12_7)*signed(FMAP_4_12);
			MULT_13(3)<=signed(DIN_13_7)*signed(FMAP_4_13);
			MULT_14(3)<=signed(DIN_14_7)*signed(FMAP_4_14);
			MULT_15(3)<=signed(DIN_15_7)*signed(FMAP_4_15);
			MULT_16(3)<=signed(DIN_16_7)*signed(FMAP_4_16);
			MULT_17(3)<=signed(DIN_17_7)*signed(FMAP_4_17);
			MULT_18(3)<=signed(DIN_18_7)*signed(FMAP_4_18);
			MULT_19(3)<=signed(DIN_19_7)*signed(FMAP_4_19);
			MULT_20(3)<=signed(DIN_20_7)*signed(FMAP_4_20);
			MULT_21(3)<=signed(DIN_21_7)*signed(FMAP_4_21);
			MULT_22(3)<=signed(DIN_22_7)*signed(FMAP_4_22);
			MULT_23(3)<=signed(DIN_23_7)*signed(FMAP_4_23);
			MULT_24(3)<=signed(DIN_24_7)*signed(FMAP_4_24);
			MULT_25(3)<=signed(DIN_25_7)*signed(FMAP_4_25);
			MULT_26(3)<=signed(DIN_26_7)*signed(FMAP_4_26);
			MULT_27(3)<=signed(DIN_27_7)*signed(FMAP_4_27);
			MULT_28(3)<=signed(DIN_28_7)*signed(FMAP_4_28);
			MULT_29(3)<=signed(DIN_29_7)*signed(FMAP_4_29);
			MULT_30(3)<=signed(DIN_30_7)*signed(FMAP_4_30);
			MULT_31(3)<=signed(DIN_31_7)*signed(FMAP_4_31);
			MULT_32(3)<=signed(DIN_32_7)*signed(FMAP_4_32);
			MULT_33(3)<=signed(DIN_33_7)*signed(FMAP_4_33);
			MULT_34(3)<=signed(DIN_34_7)*signed(FMAP_4_34);
			MULT_35(3)<=signed(DIN_35_7)*signed(FMAP_4_35);
			MULT_36(3)<=signed(DIN_36_7)*signed(FMAP_4_36);
			MULT_37(3)<=signed(DIN_37_7)*signed(FMAP_4_37);
			MULT_38(3)<=signed(DIN_38_7)*signed(FMAP_4_38);
			MULT_39(3)<=signed(DIN_39_7)*signed(FMAP_4_39);
			MULT_40(3)<=signed(DIN_40_7)*signed(FMAP_4_40);
			MULT_41(3)<=signed(DIN_41_7)*signed(FMAP_4_41);
			MULT_42(3)<=signed(DIN_42_7)*signed(FMAP_4_42);
			MULT_43(3)<=signed(DIN_43_7)*signed(FMAP_4_43);
			MULT_44(3)<=signed(DIN_44_7)*signed(FMAP_4_44);
			MULT_45(3)<=signed(DIN_45_7)*signed(FMAP_4_45);
			MULT_46(3)<=signed(DIN_46_7)*signed(FMAP_4_46);
			MULT_47(3)<=signed(DIN_47_7)*signed(FMAP_4_47);
			MULT_48(3)<=signed(DIN_48_7)*signed(FMAP_4_48);
			MULT_49(3)<=signed(DIN_49_7)*signed(FMAP_4_49);
			MULT_50(3)<=signed(DIN_50_7)*signed(FMAP_4_50);
			MULT_51(3)<=signed(DIN_51_7)*signed(FMAP_4_51);
			MULT_52(3)<=signed(DIN_52_7)*signed(FMAP_4_52);
			MULT_53(3)<=signed(DIN_53_7)*signed(FMAP_4_53);
			MULT_54(3)<=signed(DIN_54_7)*signed(FMAP_4_54);
			MULT_55(3)<=signed(DIN_55_7)*signed(FMAP_4_55);
			MULT_56(3)<=signed(DIN_56_7)*signed(FMAP_4_56);
			MULT_57(3)<=signed(DIN_57_7)*signed(FMAP_4_57);
			MULT_58(3)<=signed(DIN_58_7)*signed(FMAP_4_58);
			MULT_59(3)<=signed(DIN_59_7)*signed(FMAP_4_59);
			MULT_60(3)<=signed(DIN_60_7)*signed(FMAP_4_60);
			MULT_61(3)<=signed(DIN_61_7)*signed(FMAP_4_61);
			MULT_62(3)<=signed(DIN_62_7)*signed(FMAP_4_62);
			MULT_63(3)<=signed(DIN_63_7)*signed(FMAP_4_63);
			MULT_64(3)<=signed(DIN_64_7)*signed(FMAP_4_64);
			MULT_65(3)<=signed(DIN_65_7)*signed(FMAP_4_65);
			MULT_66(3)<=signed(DIN_66_7)*signed(FMAP_4_66);
			MULT_67(3)<=signed(DIN_67_7)*signed(FMAP_4_67);
			MULT_68(3)<=signed(DIN_68_7)*signed(FMAP_4_68);
			MULT_69(3)<=signed(DIN_69_7)*signed(FMAP_4_69);
			MULT_70(3)<=signed(DIN_70_7)*signed(FMAP_4_70);
			MULT_71(3)<=signed(DIN_71_7)*signed(FMAP_4_71);
			MULT_72(3)<=signed(DIN_72_7)*signed(FMAP_4_72);
			MULT_73(3)<=signed(DIN_73_7)*signed(FMAP_4_73);
			MULT_74(3)<=signed(DIN_74_7)*signed(FMAP_4_74);
			MULT_75(3)<=signed(DIN_75_7)*signed(FMAP_4_75);
			MULT_76(3)<=signed(DIN_76_7)*signed(FMAP_4_76);
			MULT_77(3)<=signed(DIN_77_7)*signed(FMAP_4_77);
			MULT_78(3)<=signed(DIN_78_7)*signed(FMAP_4_78);
			MULT_79(3)<=signed(DIN_79_7)*signed(FMAP_4_79);
			MULT_80(3)<=signed(DIN_80_7)*signed(FMAP_4_80);
			MULT_81(3)<=signed(DIN_81_7)*signed(FMAP_4_81);
			MULT_82(3)<=signed(DIN_82_7)*signed(FMAP_4_82);
			MULT_83(3)<=signed(DIN_83_7)*signed(FMAP_4_83);
			MULT_84(3)<=signed(DIN_84_7)*signed(FMAP_4_84);
			MULT_85(3)<=signed(DIN_85_7)*signed(FMAP_4_85);
			MULT_86(3)<=signed(DIN_86_7)*signed(FMAP_4_86);
			MULT_87(3)<=signed(DIN_87_7)*signed(FMAP_4_87);
			MULT_88(3)<=signed(DIN_88_7)*signed(FMAP_4_88);
			MULT_89(3)<=signed(DIN_89_7)*signed(FMAP_4_89);
			MULT_90(3)<=signed(DIN_90_7)*signed(FMAP_4_90);
			MULT_91(3)<=signed(DIN_91_7)*signed(FMAP_4_91);
			MULT_92(3)<=signed(DIN_92_7)*signed(FMAP_4_92);
			MULT_93(3)<=signed(DIN_93_7)*signed(FMAP_4_93);
			MULT_94(3)<=signed(DIN_94_7)*signed(FMAP_4_94);
			MULT_95(3)<=signed(DIN_95_7)*signed(FMAP_4_95);
			MULT_96(3)<=signed(DIN_96_7)*signed(FMAP_4_96);
			MULT_97(3)<=signed(DIN_97_7)*signed(FMAP_4_97);
			MULT_98(3)<=signed(DIN_98_7)*signed(FMAP_4_98);
			MULT_99(3)<=signed(DIN_99_7)*signed(FMAP_4_99);
			MULT_100(3)<=signed(DIN_100_7)*signed(FMAP_4_100);
			MULT_101(3)<=signed(DIN_101_7)*signed(FMAP_4_101);
			MULT_102(3)<=signed(DIN_102_7)*signed(FMAP_4_102);
			MULT_103(3)<=signed(DIN_103_7)*signed(FMAP_4_103);
			MULT_104(3)<=signed(DIN_104_7)*signed(FMAP_4_104);
			MULT_105(3)<=signed(DIN_105_7)*signed(FMAP_4_105);
			MULT_106(3)<=signed(DIN_106_7)*signed(FMAP_4_106);
			MULT_107(3)<=signed(DIN_107_7)*signed(FMAP_4_107);
			MULT_108(3)<=signed(DIN_108_7)*signed(FMAP_4_108);
			MULT_109(3)<=signed(DIN_109_7)*signed(FMAP_4_109);
			MULT_110(3)<=signed(DIN_110_7)*signed(FMAP_4_110);
			MULT_111(3)<=signed(DIN_111_7)*signed(FMAP_4_111);
			MULT_112(3)<=signed(DIN_112_7)*signed(FMAP_4_112);
			MULT_113(3)<=signed(DIN_113_7)*signed(FMAP_4_113);
			MULT_114(3)<=signed(DIN_114_7)*signed(FMAP_4_114);
			MULT_115(3)<=signed(DIN_115_7)*signed(FMAP_4_115);
			MULT_116(3)<=signed(DIN_116_7)*signed(FMAP_4_116);
			MULT_117(3)<=signed(DIN_117_7)*signed(FMAP_4_117);
			MULT_118(3)<=signed(DIN_118_7)*signed(FMAP_4_118);
			MULT_119(3)<=signed(DIN_119_7)*signed(FMAP_4_119);
			MULT_120(3)<=signed(DIN_120_7)*signed(FMAP_4_120);

			MULT_1(4)<=signed(DIN_1_7)*signed(FMAP_5_1);
			MULT_2(4)<=signed(DIN_2_7)*signed(FMAP_5_2);
			MULT_3(4)<=signed(DIN_3_7)*signed(FMAP_5_3);
			MULT_4(4)<=signed(DIN_4_7)*signed(FMAP_5_4);
			MULT_5(4)<=signed(DIN_5_7)*signed(FMAP_5_5);
			MULT_6(4)<=signed(DIN_6_7)*signed(FMAP_5_6);
			MULT_7(4)<=signed(DIN_7_7)*signed(FMAP_5_7);
			MULT_8(4)<=signed(DIN_8_7)*signed(FMAP_5_8);
			MULT_9(4)<=signed(DIN_9_7)*signed(FMAP_5_9);
			MULT_10(4)<=signed(DIN_10_7)*signed(FMAP_5_10);
			MULT_11(4)<=signed(DIN_11_7)*signed(FMAP_5_11);
			MULT_12(4)<=signed(DIN_12_7)*signed(FMAP_5_12);
			MULT_13(4)<=signed(DIN_13_7)*signed(FMAP_5_13);
			MULT_14(4)<=signed(DIN_14_7)*signed(FMAP_5_14);
			MULT_15(4)<=signed(DIN_15_7)*signed(FMAP_5_15);
			MULT_16(4)<=signed(DIN_16_7)*signed(FMAP_5_16);
			MULT_17(4)<=signed(DIN_17_7)*signed(FMAP_5_17);
			MULT_18(4)<=signed(DIN_18_7)*signed(FMAP_5_18);
			MULT_19(4)<=signed(DIN_19_7)*signed(FMAP_5_19);
			MULT_20(4)<=signed(DIN_20_7)*signed(FMAP_5_20);
			MULT_21(4)<=signed(DIN_21_7)*signed(FMAP_5_21);
			MULT_22(4)<=signed(DIN_22_7)*signed(FMAP_5_22);
			MULT_23(4)<=signed(DIN_23_7)*signed(FMAP_5_23);
			MULT_24(4)<=signed(DIN_24_7)*signed(FMAP_5_24);
			MULT_25(4)<=signed(DIN_25_7)*signed(FMAP_5_25);
			MULT_26(4)<=signed(DIN_26_7)*signed(FMAP_5_26);
			MULT_27(4)<=signed(DIN_27_7)*signed(FMAP_5_27);
			MULT_28(4)<=signed(DIN_28_7)*signed(FMAP_5_28);
			MULT_29(4)<=signed(DIN_29_7)*signed(FMAP_5_29);
			MULT_30(4)<=signed(DIN_30_7)*signed(FMAP_5_30);
			MULT_31(4)<=signed(DIN_31_7)*signed(FMAP_5_31);
			MULT_32(4)<=signed(DIN_32_7)*signed(FMAP_5_32);
			MULT_33(4)<=signed(DIN_33_7)*signed(FMAP_5_33);
			MULT_34(4)<=signed(DIN_34_7)*signed(FMAP_5_34);
			MULT_35(4)<=signed(DIN_35_7)*signed(FMAP_5_35);
			MULT_36(4)<=signed(DIN_36_7)*signed(FMAP_5_36);
			MULT_37(4)<=signed(DIN_37_7)*signed(FMAP_5_37);
			MULT_38(4)<=signed(DIN_38_7)*signed(FMAP_5_38);
			MULT_39(4)<=signed(DIN_39_7)*signed(FMAP_5_39);
			MULT_40(4)<=signed(DIN_40_7)*signed(FMAP_5_40);
			MULT_41(4)<=signed(DIN_41_7)*signed(FMAP_5_41);
			MULT_42(4)<=signed(DIN_42_7)*signed(FMAP_5_42);
			MULT_43(4)<=signed(DIN_43_7)*signed(FMAP_5_43);
			MULT_44(4)<=signed(DIN_44_7)*signed(FMAP_5_44);
			MULT_45(4)<=signed(DIN_45_7)*signed(FMAP_5_45);
			MULT_46(4)<=signed(DIN_46_7)*signed(FMAP_5_46);
			MULT_47(4)<=signed(DIN_47_7)*signed(FMAP_5_47);
			MULT_48(4)<=signed(DIN_48_7)*signed(FMAP_5_48);
			MULT_49(4)<=signed(DIN_49_7)*signed(FMAP_5_49);
			MULT_50(4)<=signed(DIN_50_7)*signed(FMAP_5_50);
			MULT_51(4)<=signed(DIN_51_7)*signed(FMAP_5_51);
			MULT_52(4)<=signed(DIN_52_7)*signed(FMAP_5_52);
			MULT_53(4)<=signed(DIN_53_7)*signed(FMAP_5_53);
			MULT_54(4)<=signed(DIN_54_7)*signed(FMAP_5_54);
			MULT_55(4)<=signed(DIN_55_7)*signed(FMAP_5_55);
			MULT_56(4)<=signed(DIN_56_7)*signed(FMAP_5_56);
			MULT_57(4)<=signed(DIN_57_7)*signed(FMAP_5_57);
			MULT_58(4)<=signed(DIN_58_7)*signed(FMAP_5_58);
			MULT_59(4)<=signed(DIN_59_7)*signed(FMAP_5_59);
			MULT_60(4)<=signed(DIN_60_7)*signed(FMAP_5_60);
			MULT_61(4)<=signed(DIN_61_7)*signed(FMAP_5_61);
			MULT_62(4)<=signed(DIN_62_7)*signed(FMAP_5_62);
			MULT_63(4)<=signed(DIN_63_7)*signed(FMAP_5_63);
			MULT_64(4)<=signed(DIN_64_7)*signed(FMAP_5_64);
			MULT_65(4)<=signed(DIN_65_7)*signed(FMAP_5_65);
			MULT_66(4)<=signed(DIN_66_7)*signed(FMAP_5_66);
			MULT_67(4)<=signed(DIN_67_7)*signed(FMAP_5_67);
			MULT_68(4)<=signed(DIN_68_7)*signed(FMAP_5_68);
			MULT_69(4)<=signed(DIN_69_7)*signed(FMAP_5_69);
			MULT_70(4)<=signed(DIN_70_7)*signed(FMAP_5_70);
			MULT_71(4)<=signed(DIN_71_7)*signed(FMAP_5_71);
			MULT_72(4)<=signed(DIN_72_7)*signed(FMAP_5_72);
			MULT_73(4)<=signed(DIN_73_7)*signed(FMAP_5_73);
			MULT_74(4)<=signed(DIN_74_7)*signed(FMAP_5_74);
			MULT_75(4)<=signed(DIN_75_7)*signed(FMAP_5_75);
			MULT_76(4)<=signed(DIN_76_7)*signed(FMAP_5_76);
			MULT_77(4)<=signed(DIN_77_7)*signed(FMAP_5_77);
			MULT_78(4)<=signed(DIN_78_7)*signed(FMAP_5_78);
			MULT_79(4)<=signed(DIN_79_7)*signed(FMAP_5_79);
			MULT_80(4)<=signed(DIN_80_7)*signed(FMAP_5_80);
			MULT_81(4)<=signed(DIN_81_7)*signed(FMAP_5_81);
			MULT_82(4)<=signed(DIN_82_7)*signed(FMAP_5_82);
			MULT_83(4)<=signed(DIN_83_7)*signed(FMAP_5_83);
			MULT_84(4)<=signed(DIN_84_7)*signed(FMAP_5_84);
			MULT_85(4)<=signed(DIN_85_7)*signed(FMAP_5_85);
			MULT_86(4)<=signed(DIN_86_7)*signed(FMAP_5_86);
			MULT_87(4)<=signed(DIN_87_7)*signed(FMAP_5_87);
			MULT_88(4)<=signed(DIN_88_7)*signed(FMAP_5_88);
			MULT_89(4)<=signed(DIN_89_7)*signed(FMAP_5_89);
			MULT_90(4)<=signed(DIN_90_7)*signed(FMAP_5_90);
			MULT_91(4)<=signed(DIN_91_7)*signed(FMAP_5_91);
			MULT_92(4)<=signed(DIN_92_7)*signed(FMAP_5_92);
			MULT_93(4)<=signed(DIN_93_7)*signed(FMAP_5_93);
			MULT_94(4)<=signed(DIN_94_7)*signed(FMAP_5_94);
			MULT_95(4)<=signed(DIN_95_7)*signed(FMAP_5_95);
			MULT_96(4)<=signed(DIN_96_7)*signed(FMAP_5_96);
			MULT_97(4)<=signed(DIN_97_7)*signed(FMAP_5_97);
			MULT_98(4)<=signed(DIN_98_7)*signed(FMAP_5_98);
			MULT_99(4)<=signed(DIN_99_7)*signed(FMAP_5_99);
			MULT_100(4)<=signed(DIN_100_7)*signed(FMAP_5_100);
			MULT_101(4)<=signed(DIN_101_7)*signed(FMAP_5_101);
			MULT_102(4)<=signed(DIN_102_7)*signed(FMAP_5_102);
			MULT_103(4)<=signed(DIN_103_7)*signed(FMAP_5_103);
			MULT_104(4)<=signed(DIN_104_7)*signed(FMAP_5_104);
			MULT_105(4)<=signed(DIN_105_7)*signed(FMAP_5_105);
			MULT_106(4)<=signed(DIN_106_7)*signed(FMAP_5_106);
			MULT_107(4)<=signed(DIN_107_7)*signed(FMAP_5_107);
			MULT_108(4)<=signed(DIN_108_7)*signed(FMAP_5_108);
			MULT_109(4)<=signed(DIN_109_7)*signed(FMAP_5_109);
			MULT_110(4)<=signed(DIN_110_7)*signed(FMAP_5_110);
			MULT_111(4)<=signed(DIN_111_7)*signed(FMAP_5_111);
			MULT_112(4)<=signed(DIN_112_7)*signed(FMAP_5_112);
			MULT_113(4)<=signed(DIN_113_7)*signed(FMAP_5_113);
			MULT_114(4)<=signed(DIN_114_7)*signed(FMAP_5_114);
			MULT_115(4)<=signed(DIN_115_7)*signed(FMAP_5_115);
			MULT_116(4)<=signed(DIN_116_7)*signed(FMAP_5_116);
			MULT_117(4)<=signed(DIN_117_7)*signed(FMAP_5_117);
			MULT_118(4)<=signed(DIN_118_7)*signed(FMAP_5_118);
			MULT_119(4)<=signed(DIN_119_7)*signed(FMAP_5_119);
			MULT_120(4)<=signed(DIN_120_7)*signed(FMAP_5_120);

			MULT_1(5)<=signed(DIN_1_7)*signed(FMAP_6_1);
			MULT_2(5)<=signed(DIN_2_7)*signed(FMAP_6_2);
			MULT_3(5)<=signed(DIN_3_7)*signed(FMAP_6_3);
			MULT_4(5)<=signed(DIN_4_7)*signed(FMAP_6_4);
			MULT_5(5)<=signed(DIN_5_7)*signed(FMAP_6_5);
			MULT_6(5)<=signed(DIN_6_7)*signed(FMAP_6_6);
			MULT_7(5)<=signed(DIN_7_7)*signed(FMAP_6_7);
			MULT_8(5)<=signed(DIN_8_7)*signed(FMAP_6_8);
			MULT_9(5)<=signed(DIN_9_7)*signed(FMAP_6_9);
			MULT_10(5)<=signed(DIN_10_7)*signed(FMAP_6_10);
			MULT_11(5)<=signed(DIN_11_7)*signed(FMAP_6_11);
			MULT_12(5)<=signed(DIN_12_7)*signed(FMAP_6_12);
			MULT_13(5)<=signed(DIN_13_7)*signed(FMAP_6_13);
			MULT_14(5)<=signed(DIN_14_7)*signed(FMAP_6_14);
			MULT_15(5)<=signed(DIN_15_7)*signed(FMAP_6_15);
			MULT_16(5)<=signed(DIN_16_7)*signed(FMAP_6_16);
			MULT_17(5)<=signed(DIN_17_7)*signed(FMAP_6_17);
			MULT_18(5)<=signed(DIN_18_7)*signed(FMAP_6_18);
			MULT_19(5)<=signed(DIN_19_7)*signed(FMAP_6_19);
			MULT_20(5)<=signed(DIN_20_7)*signed(FMAP_6_20);
			MULT_21(5)<=signed(DIN_21_7)*signed(FMAP_6_21);
			MULT_22(5)<=signed(DIN_22_7)*signed(FMAP_6_22);
			MULT_23(5)<=signed(DIN_23_7)*signed(FMAP_6_23);
			MULT_24(5)<=signed(DIN_24_7)*signed(FMAP_6_24);
			MULT_25(5)<=signed(DIN_25_7)*signed(FMAP_6_25);
			MULT_26(5)<=signed(DIN_26_7)*signed(FMAP_6_26);
			MULT_27(5)<=signed(DIN_27_7)*signed(FMAP_6_27);
			MULT_28(5)<=signed(DIN_28_7)*signed(FMAP_6_28);
			MULT_29(5)<=signed(DIN_29_7)*signed(FMAP_6_29);
			MULT_30(5)<=signed(DIN_30_7)*signed(FMAP_6_30);
			MULT_31(5)<=signed(DIN_31_7)*signed(FMAP_6_31);
			MULT_32(5)<=signed(DIN_32_7)*signed(FMAP_6_32);
			MULT_33(5)<=signed(DIN_33_7)*signed(FMAP_6_33);
			MULT_34(5)<=signed(DIN_34_7)*signed(FMAP_6_34);
			MULT_35(5)<=signed(DIN_35_7)*signed(FMAP_6_35);
			MULT_36(5)<=signed(DIN_36_7)*signed(FMAP_6_36);
			MULT_37(5)<=signed(DIN_37_7)*signed(FMAP_6_37);
			MULT_38(5)<=signed(DIN_38_7)*signed(FMAP_6_38);
			MULT_39(5)<=signed(DIN_39_7)*signed(FMAP_6_39);
			MULT_40(5)<=signed(DIN_40_7)*signed(FMAP_6_40);
			MULT_41(5)<=signed(DIN_41_7)*signed(FMAP_6_41);
			MULT_42(5)<=signed(DIN_42_7)*signed(FMAP_6_42);
			MULT_43(5)<=signed(DIN_43_7)*signed(FMAP_6_43);
			MULT_44(5)<=signed(DIN_44_7)*signed(FMAP_6_44);
			MULT_45(5)<=signed(DIN_45_7)*signed(FMAP_6_45);
			MULT_46(5)<=signed(DIN_46_7)*signed(FMAP_6_46);
			MULT_47(5)<=signed(DIN_47_7)*signed(FMAP_6_47);
			MULT_48(5)<=signed(DIN_48_7)*signed(FMAP_6_48);
			MULT_49(5)<=signed(DIN_49_7)*signed(FMAP_6_49);
			MULT_50(5)<=signed(DIN_50_7)*signed(FMAP_6_50);
			MULT_51(5)<=signed(DIN_51_7)*signed(FMAP_6_51);
			MULT_52(5)<=signed(DIN_52_7)*signed(FMAP_6_52);
			MULT_53(5)<=signed(DIN_53_7)*signed(FMAP_6_53);
			MULT_54(5)<=signed(DIN_54_7)*signed(FMAP_6_54);
			MULT_55(5)<=signed(DIN_55_7)*signed(FMAP_6_55);
			MULT_56(5)<=signed(DIN_56_7)*signed(FMAP_6_56);
			MULT_57(5)<=signed(DIN_57_7)*signed(FMAP_6_57);
			MULT_58(5)<=signed(DIN_58_7)*signed(FMAP_6_58);
			MULT_59(5)<=signed(DIN_59_7)*signed(FMAP_6_59);
			MULT_60(5)<=signed(DIN_60_7)*signed(FMAP_6_60);
			MULT_61(5)<=signed(DIN_61_7)*signed(FMAP_6_61);
			MULT_62(5)<=signed(DIN_62_7)*signed(FMAP_6_62);
			MULT_63(5)<=signed(DIN_63_7)*signed(FMAP_6_63);
			MULT_64(5)<=signed(DIN_64_7)*signed(FMAP_6_64);
			MULT_65(5)<=signed(DIN_65_7)*signed(FMAP_6_65);
			MULT_66(5)<=signed(DIN_66_7)*signed(FMAP_6_66);
			MULT_67(5)<=signed(DIN_67_7)*signed(FMAP_6_67);
			MULT_68(5)<=signed(DIN_68_7)*signed(FMAP_6_68);
			MULT_69(5)<=signed(DIN_69_7)*signed(FMAP_6_69);
			MULT_70(5)<=signed(DIN_70_7)*signed(FMAP_6_70);
			MULT_71(5)<=signed(DIN_71_7)*signed(FMAP_6_71);
			MULT_72(5)<=signed(DIN_72_7)*signed(FMAP_6_72);
			MULT_73(5)<=signed(DIN_73_7)*signed(FMAP_6_73);
			MULT_74(5)<=signed(DIN_74_7)*signed(FMAP_6_74);
			MULT_75(5)<=signed(DIN_75_7)*signed(FMAP_6_75);
			MULT_76(5)<=signed(DIN_76_7)*signed(FMAP_6_76);
			MULT_77(5)<=signed(DIN_77_7)*signed(FMAP_6_77);
			MULT_78(5)<=signed(DIN_78_7)*signed(FMAP_6_78);
			MULT_79(5)<=signed(DIN_79_7)*signed(FMAP_6_79);
			MULT_80(5)<=signed(DIN_80_7)*signed(FMAP_6_80);
			MULT_81(5)<=signed(DIN_81_7)*signed(FMAP_6_81);
			MULT_82(5)<=signed(DIN_82_7)*signed(FMAP_6_82);
			MULT_83(5)<=signed(DIN_83_7)*signed(FMAP_6_83);
			MULT_84(5)<=signed(DIN_84_7)*signed(FMAP_6_84);
			MULT_85(5)<=signed(DIN_85_7)*signed(FMAP_6_85);
			MULT_86(5)<=signed(DIN_86_7)*signed(FMAP_6_86);
			MULT_87(5)<=signed(DIN_87_7)*signed(FMAP_6_87);
			MULT_88(5)<=signed(DIN_88_7)*signed(FMAP_6_88);
			MULT_89(5)<=signed(DIN_89_7)*signed(FMAP_6_89);
			MULT_90(5)<=signed(DIN_90_7)*signed(FMAP_6_90);
			MULT_91(5)<=signed(DIN_91_7)*signed(FMAP_6_91);
			MULT_92(5)<=signed(DIN_92_7)*signed(FMAP_6_92);
			MULT_93(5)<=signed(DIN_93_7)*signed(FMAP_6_93);
			MULT_94(5)<=signed(DIN_94_7)*signed(FMAP_6_94);
			MULT_95(5)<=signed(DIN_95_7)*signed(FMAP_6_95);
			MULT_96(5)<=signed(DIN_96_7)*signed(FMAP_6_96);
			MULT_97(5)<=signed(DIN_97_7)*signed(FMAP_6_97);
			MULT_98(5)<=signed(DIN_98_7)*signed(FMAP_6_98);
			MULT_99(5)<=signed(DIN_99_7)*signed(FMAP_6_99);
			MULT_100(5)<=signed(DIN_100_7)*signed(FMAP_6_100);
			MULT_101(5)<=signed(DIN_101_7)*signed(FMAP_6_101);
			MULT_102(5)<=signed(DIN_102_7)*signed(FMAP_6_102);
			MULT_103(5)<=signed(DIN_103_7)*signed(FMAP_6_103);
			MULT_104(5)<=signed(DIN_104_7)*signed(FMAP_6_104);
			MULT_105(5)<=signed(DIN_105_7)*signed(FMAP_6_105);
			MULT_106(5)<=signed(DIN_106_7)*signed(FMAP_6_106);
			MULT_107(5)<=signed(DIN_107_7)*signed(FMAP_6_107);
			MULT_108(5)<=signed(DIN_108_7)*signed(FMAP_6_108);
			MULT_109(5)<=signed(DIN_109_7)*signed(FMAP_6_109);
			MULT_110(5)<=signed(DIN_110_7)*signed(FMAP_6_110);
			MULT_111(5)<=signed(DIN_111_7)*signed(FMAP_6_111);
			MULT_112(5)<=signed(DIN_112_7)*signed(FMAP_6_112);
			MULT_113(5)<=signed(DIN_113_7)*signed(FMAP_6_113);
			MULT_114(5)<=signed(DIN_114_7)*signed(FMAP_6_114);
			MULT_115(5)<=signed(DIN_115_7)*signed(FMAP_6_115);
			MULT_116(5)<=signed(DIN_116_7)*signed(FMAP_6_116);
			MULT_117(5)<=signed(DIN_117_7)*signed(FMAP_6_117);
			MULT_118(5)<=signed(DIN_118_7)*signed(FMAP_6_118);
			MULT_119(5)<=signed(DIN_119_7)*signed(FMAP_6_119);
			MULT_120(5)<=signed(DIN_120_7)*signed(FMAP_6_120);

			MULT_1(6)<=signed(DIN_1_7)*signed(FMAP_7_1);
			MULT_2(6)<=signed(DIN_2_7)*signed(FMAP_7_2);
			MULT_3(6)<=signed(DIN_3_7)*signed(FMAP_7_3);
			MULT_4(6)<=signed(DIN_4_7)*signed(FMAP_7_4);
			MULT_5(6)<=signed(DIN_5_7)*signed(FMAP_7_5);
			MULT_6(6)<=signed(DIN_6_7)*signed(FMAP_7_6);
			MULT_7(6)<=signed(DIN_7_7)*signed(FMAP_7_7);
			MULT_8(6)<=signed(DIN_8_7)*signed(FMAP_7_8);
			MULT_9(6)<=signed(DIN_9_7)*signed(FMAP_7_9);
			MULT_10(6)<=signed(DIN_10_7)*signed(FMAP_7_10);
			MULT_11(6)<=signed(DIN_11_7)*signed(FMAP_7_11);
			MULT_12(6)<=signed(DIN_12_7)*signed(FMAP_7_12);
			MULT_13(6)<=signed(DIN_13_7)*signed(FMAP_7_13);
			MULT_14(6)<=signed(DIN_14_7)*signed(FMAP_7_14);
			MULT_15(6)<=signed(DIN_15_7)*signed(FMAP_7_15);
			MULT_16(6)<=signed(DIN_16_7)*signed(FMAP_7_16);
			MULT_17(6)<=signed(DIN_17_7)*signed(FMAP_7_17);
			MULT_18(6)<=signed(DIN_18_7)*signed(FMAP_7_18);
			MULT_19(6)<=signed(DIN_19_7)*signed(FMAP_7_19);
			MULT_20(6)<=signed(DIN_20_7)*signed(FMAP_7_20);
			MULT_21(6)<=signed(DIN_21_7)*signed(FMAP_7_21);
			MULT_22(6)<=signed(DIN_22_7)*signed(FMAP_7_22);
			MULT_23(6)<=signed(DIN_23_7)*signed(FMAP_7_23);
			MULT_24(6)<=signed(DIN_24_7)*signed(FMAP_7_24);
			MULT_25(6)<=signed(DIN_25_7)*signed(FMAP_7_25);
			MULT_26(6)<=signed(DIN_26_7)*signed(FMAP_7_26);
			MULT_27(6)<=signed(DIN_27_7)*signed(FMAP_7_27);
			MULT_28(6)<=signed(DIN_28_7)*signed(FMAP_7_28);
			MULT_29(6)<=signed(DIN_29_7)*signed(FMAP_7_29);
			MULT_30(6)<=signed(DIN_30_7)*signed(FMAP_7_30);
			MULT_31(6)<=signed(DIN_31_7)*signed(FMAP_7_31);
			MULT_32(6)<=signed(DIN_32_7)*signed(FMAP_7_32);
			MULT_33(6)<=signed(DIN_33_7)*signed(FMAP_7_33);
			MULT_34(6)<=signed(DIN_34_7)*signed(FMAP_7_34);
			MULT_35(6)<=signed(DIN_35_7)*signed(FMAP_7_35);
			MULT_36(6)<=signed(DIN_36_7)*signed(FMAP_7_36);
			MULT_37(6)<=signed(DIN_37_7)*signed(FMAP_7_37);
			MULT_38(6)<=signed(DIN_38_7)*signed(FMAP_7_38);
			MULT_39(6)<=signed(DIN_39_7)*signed(FMAP_7_39);
			MULT_40(6)<=signed(DIN_40_7)*signed(FMAP_7_40);
			MULT_41(6)<=signed(DIN_41_7)*signed(FMAP_7_41);
			MULT_42(6)<=signed(DIN_42_7)*signed(FMAP_7_42);
			MULT_43(6)<=signed(DIN_43_7)*signed(FMAP_7_43);
			MULT_44(6)<=signed(DIN_44_7)*signed(FMAP_7_44);
			MULT_45(6)<=signed(DIN_45_7)*signed(FMAP_7_45);
			MULT_46(6)<=signed(DIN_46_7)*signed(FMAP_7_46);
			MULT_47(6)<=signed(DIN_47_7)*signed(FMAP_7_47);
			MULT_48(6)<=signed(DIN_48_7)*signed(FMAP_7_48);
			MULT_49(6)<=signed(DIN_49_7)*signed(FMAP_7_49);
			MULT_50(6)<=signed(DIN_50_7)*signed(FMAP_7_50);
			MULT_51(6)<=signed(DIN_51_7)*signed(FMAP_7_51);
			MULT_52(6)<=signed(DIN_52_7)*signed(FMAP_7_52);
			MULT_53(6)<=signed(DIN_53_7)*signed(FMAP_7_53);
			MULT_54(6)<=signed(DIN_54_7)*signed(FMAP_7_54);
			MULT_55(6)<=signed(DIN_55_7)*signed(FMAP_7_55);
			MULT_56(6)<=signed(DIN_56_7)*signed(FMAP_7_56);
			MULT_57(6)<=signed(DIN_57_7)*signed(FMAP_7_57);
			MULT_58(6)<=signed(DIN_58_7)*signed(FMAP_7_58);
			MULT_59(6)<=signed(DIN_59_7)*signed(FMAP_7_59);
			MULT_60(6)<=signed(DIN_60_7)*signed(FMAP_7_60);
			MULT_61(6)<=signed(DIN_61_7)*signed(FMAP_7_61);
			MULT_62(6)<=signed(DIN_62_7)*signed(FMAP_7_62);
			MULT_63(6)<=signed(DIN_63_7)*signed(FMAP_7_63);
			MULT_64(6)<=signed(DIN_64_7)*signed(FMAP_7_64);
			MULT_65(6)<=signed(DIN_65_7)*signed(FMAP_7_65);
			MULT_66(6)<=signed(DIN_66_7)*signed(FMAP_7_66);
			MULT_67(6)<=signed(DIN_67_7)*signed(FMAP_7_67);
			MULT_68(6)<=signed(DIN_68_7)*signed(FMAP_7_68);
			MULT_69(6)<=signed(DIN_69_7)*signed(FMAP_7_69);
			MULT_70(6)<=signed(DIN_70_7)*signed(FMAP_7_70);
			MULT_71(6)<=signed(DIN_71_7)*signed(FMAP_7_71);
			MULT_72(6)<=signed(DIN_72_7)*signed(FMAP_7_72);
			MULT_73(6)<=signed(DIN_73_7)*signed(FMAP_7_73);
			MULT_74(6)<=signed(DIN_74_7)*signed(FMAP_7_74);
			MULT_75(6)<=signed(DIN_75_7)*signed(FMAP_7_75);
			MULT_76(6)<=signed(DIN_76_7)*signed(FMAP_7_76);
			MULT_77(6)<=signed(DIN_77_7)*signed(FMAP_7_77);
			MULT_78(6)<=signed(DIN_78_7)*signed(FMAP_7_78);
			MULT_79(6)<=signed(DIN_79_7)*signed(FMAP_7_79);
			MULT_80(6)<=signed(DIN_80_7)*signed(FMAP_7_80);
			MULT_81(6)<=signed(DIN_81_7)*signed(FMAP_7_81);
			MULT_82(6)<=signed(DIN_82_7)*signed(FMAP_7_82);
			MULT_83(6)<=signed(DIN_83_7)*signed(FMAP_7_83);
			MULT_84(6)<=signed(DIN_84_7)*signed(FMAP_7_84);
			MULT_85(6)<=signed(DIN_85_7)*signed(FMAP_7_85);
			MULT_86(6)<=signed(DIN_86_7)*signed(FMAP_7_86);
			MULT_87(6)<=signed(DIN_87_7)*signed(FMAP_7_87);
			MULT_88(6)<=signed(DIN_88_7)*signed(FMAP_7_88);
			MULT_89(6)<=signed(DIN_89_7)*signed(FMAP_7_89);
			MULT_90(6)<=signed(DIN_90_7)*signed(FMAP_7_90);
			MULT_91(6)<=signed(DIN_91_7)*signed(FMAP_7_91);
			MULT_92(6)<=signed(DIN_92_7)*signed(FMAP_7_92);
			MULT_93(6)<=signed(DIN_93_7)*signed(FMAP_7_93);
			MULT_94(6)<=signed(DIN_94_7)*signed(FMAP_7_94);
			MULT_95(6)<=signed(DIN_95_7)*signed(FMAP_7_95);
			MULT_96(6)<=signed(DIN_96_7)*signed(FMAP_7_96);
			MULT_97(6)<=signed(DIN_97_7)*signed(FMAP_7_97);
			MULT_98(6)<=signed(DIN_98_7)*signed(FMAP_7_98);
			MULT_99(6)<=signed(DIN_99_7)*signed(FMAP_7_99);
			MULT_100(6)<=signed(DIN_100_7)*signed(FMAP_7_100);
			MULT_101(6)<=signed(DIN_101_7)*signed(FMAP_7_101);
			MULT_102(6)<=signed(DIN_102_7)*signed(FMAP_7_102);
			MULT_103(6)<=signed(DIN_103_7)*signed(FMAP_7_103);
			MULT_104(6)<=signed(DIN_104_7)*signed(FMAP_7_104);
			MULT_105(6)<=signed(DIN_105_7)*signed(FMAP_7_105);
			MULT_106(6)<=signed(DIN_106_7)*signed(FMAP_7_106);
			MULT_107(6)<=signed(DIN_107_7)*signed(FMAP_7_107);
			MULT_108(6)<=signed(DIN_108_7)*signed(FMAP_7_108);
			MULT_109(6)<=signed(DIN_109_7)*signed(FMAP_7_109);
			MULT_110(6)<=signed(DIN_110_7)*signed(FMAP_7_110);
			MULT_111(6)<=signed(DIN_111_7)*signed(FMAP_7_111);
			MULT_112(6)<=signed(DIN_112_7)*signed(FMAP_7_112);
			MULT_113(6)<=signed(DIN_113_7)*signed(FMAP_7_113);
			MULT_114(6)<=signed(DIN_114_7)*signed(FMAP_7_114);
			MULT_115(6)<=signed(DIN_115_7)*signed(FMAP_7_115);
			MULT_116(6)<=signed(DIN_116_7)*signed(FMAP_7_116);
			MULT_117(6)<=signed(DIN_117_7)*signed(FMAP_7_117);
			MULT_118(6)<=signed(DIN_118_7)*signed(FMAP_7_118);
			MULT_119(6)<=signed(DIN_119_7)*signed(FMAP_7_119);
			MULT_120(6)<=signed(DIN_120_7)*signed(FMAP_7_120);

			MULT_1(7)<=signed(DIN_1_7)*signed(FMAP_8_1);
			MULT_2(7)<=signed(DIN_2_7)*signed(FMAP_8_2);
			MULT_3(7)<=signed(DIN_3_7)*signed(FMAP_8_3);
			MULT_4(7)<=signed(DIN_4_7)*signed(FMAP_8_4);
			MULT_5(7)<=signed(DIN_5_7)*signed(FMAP_8_5);
			MULT_6(7)<=signed(DIN_6_7)*signed(FMAP_8_6);
			MULT_7(7)<=signed(DIN_7_7)*signed(FMAP_8_7);
			MULT_8(7)<=signed(DIN_8_7)*signed(FMAP_8_8);
			MULT_9(7)<=signed(DIN_9_7)*signed(FMAP_8_9);
			MULT_10(7)<=signed(DIN_10_7)*signed(FMAP_8_10);
			MULT_11(7)<=signed(DIN_11_7)*signed(FMAP_8_11);
			MULT_12(7)<=signed(DIN_12_7)*signed(FMAP_8_12);
			MULT_13(7)<=signed(DIN_13_7)*signed(FMAP_8_13);
			MULT_14(7)<=signed(DIN_14_7)*signed(FMAP_8_14);
			MULT_15(7)<=signed(DIN_15_7)*signed(FMAP_8_15);
			MULT_16(7)<=signed(DIN_16_7)*signed(FMAP_8_16);
			MULT_17(7)<=signed(DIN_17_7)*signed(FMAP_8_17);
			MULT_18(7)<=signed(DIN_18_7)*signed(FMAP_8_18);
			MULT_19(7)<=signed(DIN_19_7)*signed(FMAP_8_19);
			MULT_20(7)<=signed(DIN_20_7)*signed(FMAP_8_20);
			MULT_21(7)<=signed(DIN_21_7)*signed(FMAP_8_21);
			MULT_22(7)<=signed(DIN_22_7)*signed(FMAP_8_22);
			MULT_23(7)<=signed(DIN_23_7)*signed(FMAP_8_23);
			MULT_24(7)<=signed(DIN_24_7)*signed(FMAP_8_24);
			MULT_25(7)<=signed(DIN_25_7)*signed(FMAP_8_25);
			MULT_26(7)<=signed(DIN_26_7)*signed(FMAP_8_26);
			MULT_27(7)<=signed(DIN_27_7)*signed(FMAP_8_27);
			MULT_28(7)<=signed(DIN_28_7)*signed(FMAP_8_28);
			MULT_29(7)<=signed(DIN_29_7)*signed(FMAP_8_29);
			MULT_30(7)<=signed(DIN_30_7)*signed(FMAP_8_30);
			MULT_31(7)<=signed(DIN_31_7)*signed(FMAP_8_31);
			MULT_32(7)<=signed(DIN_32_7)*signed(FMAP_8_32);
			MULT_33(7)<=signed(DIN_33_7)*signed(FMAP_8_33);
			MULT_34(7)<=signed(DIN_34_7)*signed(FMAP_8_34);
			MULT_35(7)<=signed(DIN_35_7)*signed(FMAP_8_35);
			MULT_36(7)<=signed(DIN_36_7)*signed(FMAP_8_36);
			MULT_37(7)<=signed(DIN_37_7)*signed(FMAP_8_37);
			MULT_38(7)<=signed(DIN_38_7)*signed(FMAP_8_38);
			MULT_39(7)<=signed(DIN_39_7)*signed(FMAP_8_39);
			MULT_40(7)<=signed(DIN_40_7)*signed(FMAP_8_40);
			MULT_41(7)<=signed(DIN_41_7)*signed(FMAP_8_41);
			MULT_42(7)<=signed(DIN_42_7)*signed(FMAP_8_42);
			MULT_43(7)<=signed(DIN_43_7)*signed(FMAP_8_43);
			MULT_44(7)<=signed(DIN_44_7)*signed(FMAP_8_44);
			MULT_45(7)<=signed(DIN_45_7)*signed(FMAP_8_45);
			MULT_46(7)<=signed(DIN_46_7)*signed(FMAP_8_46);
			MULT_47(7)<=signed(DIN_47_7)*signed(FMAP_8_47);
			MULT_48(7)<=signed(DIN_48_7)*signed(FMAP_8_48);
			MULT_49(7)<=signed(DIN_49_7)*signed(FMAP_8_49);
			MULT_50(7)<=signed(DIN_50_7)*signed(FMAP_8_50);
			MULT_51(7)<=signed(DIN_51_7)*signed(FMAP_8_51);
			MULT_52(7)<=signed(DIN_52_7)*signed(FMAP_8_52);
			MULT_53(7)<=signed(DIN_53_7)*signed(FMAP_8_53);
			MULT_54(7)<=signed(DIN_54_7)*signed(FMAP_8_54);
			MULT_55(7)<=signed(DIN_55_7)*signed(FMAP_8_55);
			MULT_56(7)<=signed(DIN_56_7)*signed(FMAP_8_56);
			MULT_57(7)<=signed(DIN_57_7)*signed(FMAP_8_57);
			MULT_58(7)<=signed(DIN_58_7)*signed(FMAP_8_58);
			MULT_59(7)<=signed(DIN_59_7)*signed(FMAP_8_59);
			MULT_60(7)<=signed(DIN_60_7)*signed(FMAP_8_60);
			MULT_61(7)<=signed(DIN_61_7)*signed(FMAP_8_61);
			MULT_62(7)<=signed(DIN_62_7)*signed(FMAP_8_62);
			MULT_63(7)<=signed(DIN_63_7)*signed(FMAP_8_63);
			MULT_64(7)<=signed(DIN_64_7)*signed(FMAP_8_64);
			MULT_65(7)<=signed(DIN_65_7)*signed(FMAP_8_65);
			MULT_66(7)<=signed(DIN_66_7)*signed(FMAP_8_66);
			MULT_67(7)<=signed(DIN_67_7)*signed(FMAP_8_67);
			MULT_68(7)<=signed(DIN_68_7)*signed(FMAP_8_68);
			MULT_69(7)<=signed(DIN_69_7)*signed(FMAP_8_69);
			MULT_70(7)<=signed(DIN_70_7)*signed(FMAP_8_70);
			MULT_71(7)<=signed(DIN_71_7)*signed(FMAP_8_71);
			MULT_72(7)<=signed(DIN_72_7)*signed(FMAP_8_72);
			MULT_73(7)<=signed(DIN_73_7)*signed(FMAP_8_73);
			MULT_74(7)<=signed(DIN_74_7)*signed(FMAP_8_74);
			MULT_75(7)<=signed(DIN_75_7)*signed(FMAP_8_75);
			MULT_76(7)<=signed(DIN_76_7)*signed(FMAP_8_76);
			MULT_77(7)<=signed(DIN_77_7)*signed(FMAP_8_77);
			MULT_78(7)<=signed(DIN_78_7)*signed(FMAP_8_78);
			MULT_79(7)<=signed(DIN_79_7)*signed(FMAP_8_79);
			MULT_80(7)<=signed(DIN_80_7)*signed(FMAP_8_80);
			MULT_81(7)<=signed(DIN_81_7)*signed(FMAP_8_81);
			MULT_82(7)<=signed(DIN_82_7)*signed(FMAP_8_82);
			MULT_83(7)<=signed(DIN_83_7)*signed(FMAP_8_83);
			MULT_84(7)<=signed(DIN_84_7)*signed(FMAP_8_84);
			MULT_85(7)<=signed(DIN_85_7)*signed(FMAP_8_85);
			MULT_86(7)<=signed(DIN_86_7)*signed(FMAP_8_86);
			MULT_87(7)<=signed(DIN_87_7)*signed(FMAP_8_87);
			MULT_88(7)<=signed(DIN_88_7)*signed(FMAP_8_88);
			MULT_89(7)<=signed(DIN_89_7)*signed(FMAP_8_89);
			MULT_90(7)<=signed(DIN_90_7)*signed(FMAP_8_90);
			MULT_91(7)<=signed(DIN_91_7)*signed(FMAP_8_91);
			MULT_92(7)<=signed(DIN_92_7)*signed(FMAP_8_92);
			MULT_93(7)<=signed(DIN_93_7)*signed(FMAP_8_93);
			MULT_94(7)<=signed(DIN_94_7)*signed(FMAP_8_94);
			MULT_95(7)<=signed(DIN_95_7)*signed(FMAP_8_95);
			MULT_96(7)<=signed(DIN_96_7)*signed(FMAP_8_96);
			MULT_97(7)<=signed(DIN_97_7)*signed(FMAP_8_97);
			MULT_98(7)<=signed(DIN_98_7)*signed(FMAP_8_98);
			MULT_99(7)<=signed(DIN_99_7)*signed(FMAP_8_99);
			MULT_100(7)<=signed(DIN_100_7)*signed(FMAP_8_100);
			MULT_101(7)<=signed(DIN_101_7)*signed(FMAP_8_101);
			MULT_102(7)<=signed(DIN_102_7)*signed(FMAP_8_102);
			MULT_103(7)<=signed(DIN_103_7)*signed(FMAP_8_103);
			MULT_104(7)<=signed(DIN_104_7)*signed(FMAP_8_104);
			MULT_105(7)<=signed(DIN_105_7)*signed(FMAP_8_105);
			MULT_106(7)<=signed(DIN_106_7)*signed(FMAP_8_106);
			MULT_107(7)<=signed(DIN_107_7)*signed(FMAP_8_107);
			MULT_108(7)<=signed(DIN_108_7)*signed(FMAP_8_108);
			MULT_109(7)<=signed(DIN_109_7)*signed(FMAP_8_109);
			MULT_110(7)<=signed(DIN_110_7)*signed(FMAP_8_110);
			MULT_111(7)<=signed(DIN_111_7)*signed(FMAP_8_111);
			MULT_112(7)<=signed(DIN_112_7)*signed(FMAP_8_112);
			MULT_113(7)<=signed(DIN_113_7)*signed(FMAP_8_113);
			MULT_114(7)<=signed(DIN_114_7)*signed(FMAP_8_114);
			MULT_115(7)<=signed(DIN_115_7)*signed(FMAP_8_115);
			MULT_116(7)<=signed(DIN_116_7)*signed(FMAP_8_116);
			MULT_117(7)<=signed(DIN_117_7)*signed(FMAP_8_117);
			MULT_118(7)<=signed(DIN_118_7)*signed(FMAP_8_118);
			MULT_119(7)<=signed(DIN_119_7)*signed(FMAP_8_119);
			MULT_120(7)<=signed(DIN_120_7)*signed(FMAP_8_120);

			MULT_1(8)<=signed(DIN_1_7)*signed(FMAP_9_1);
			MULT_2(8)<=signed(DIN_2_7)*signed(FMAP_9_2);
			MULT_3(8)<=signed(DIN_3_7)*signed(FMAP_9_3);
			MULT_4(8)<=signed(DIN_4_7)*signed(FMAP_9_4);
			MULT_5(8)<=signed(DIN_5_7)*signed(FMAP_9_5);
			MULT_6(8)<=signed(DIN_6_7)*signed(FMAP_9_6);
			MULT_7(8)<=signed(DIN_7_7)*signed(FMAP_9_7);
			MULT_8(8)<=signed(DIN_8_7)*signed(FMAP_9_8);
			MULT_9(8)<=signed(DIN_9_7)*signed(FMAP_9_9);
			MULT_10(8)<=signed(DIN_10_7)*signed(FMAP_9_10);
			MULT_11(8)<=signed(DIN_11_7)*signed(FMAP_9_11);
			MULT_12(8)<=signed(DIN_12_7)*signed(FMAP_9_12);
			MULT_13(8)<=signed(DIN_13_7)*signed(FMAP_9_13);
			MULT_14(8)<=signed(DIN_14_7)*signed(FMAP_9_14);
			MULT_15(8)<=signed(DIN_15_7)*signed(FMAP_9_15);
			MULT_16(8)<=signed(DIN_16_7)*signed(FMAP_9_16);
			MULT_17(8)<=signed(DIN_17_7)*signed(FMAP_9_17);
			MULT_18(8)<=signed(DIN_18_7)*signed(FMAP_9_18);
			MULT_19(8)<=signed(DIN_19_7)*signed(FMAP_9_19);
			MULT_20(8)<=signed(DIN_20_7)*signed(FMAP_9_20);
			MULT_21(8)<=signed(DIN_21_7)*signed(FMAP_9_21);
			MULT_22(8)<=signed(DIN_22_7)*signed(FMAP_9_22);
			MULT_23(8)<=signed(DIN_23_7)*signed(FMAP_9_23);
			MULT_24(8)<=signed(DIN_24_7)*signed(FMAP_9_24);
			MULT_25(8)<=signed(DIN_25_7)*signed(FMAP_9_25);
			MULT_26(8)<=signed(DIN_26_7)*signed(FMAP_9_26);
			MULT_27(8)<=signed(DIN_27_7)*signed(FMAP_9_27);
			MULT_28(8)<=signed(DIN_28_7)*signed(FMAP_9_28);
			MULT_29(8)<=signed(DIN_29_7)*signed(FMAP_9_29);
			MULT_30(8)<=signed(DIN_30_7)*signed(FMAP_9_30);
			MULT_31(8)<=signed(DIN_31_7)*signed(FMAP_9_31);
			MULT_32(8)<=signed(DIN_32_7)*signed(FMAP_9_32);
			MULT_33(8)<=signed(DIN_33_7)*signed(FMAP_9_33);
			MULT_34(8)<=signed(DIN_34_7)*signed(FMAP_9_34);
			MULT_35(8)<=signed(DIN_35_7)*signed(FMAP_9_35);
			MULT_36(8)<=signed(DIN_36_7)*signed(FMAP_9_36);
			MULT_37(8)<=signed(DIN_37_7)*signed(FMAP_9_37);
			MULT_38(8)<=signed(DIN_38_7)*signed(FMAP_9_38);
			MULT_39(8)<=signed(DIN_39_7)*signed(FMAP_9_39);
			MULT_40(8)<=signed(DIN_40_7)*signed(FMAP_9_40);
			MULT_41(8)<=signed(DIN_41_7)*signed(FMAP_9_41);
			MULT_42(8)<=signed(DIN_42_7)*signed(FMAP_9_42);
			MULT_43(8)<=signed(DIN_43_7)*signed(FMAP_9_43);
			MULT_44(8)<=signed(DIN_44_7)*signed(FMAP_9_44);
			MULT_45(8)<=signed(DIN_45_7)*signed(FMAP_9_45);
			MULT_46(8)<=signed(DIN_46_7)*signed(FMAP_9_46);
			MULT_47(8)<=signed(DIN_47_7)*signed(FMAP_9_47);
			MULT_48(8)<=signed(DIN_48_7)*signed(FMAP_9_48);
			MULT_49(8)<=signed(DIN_49_7)*signed(FMAP_9_49);
			MULT_50(8)<=signed(DIN_50_7)*signed(FMAP_9_50);
			MULT_51(8)<=signed(DIN_51_7)*signed(FMAP_9_51);
			MULT_52(8)<=signed(DIN_52_7)*signed(FMAP_9_52);
			MULT_53(8)<=signed(DIN_53_7)*signed(FMAP_9_53);
			MULT_54(8)<=signed(DIN_54_7)*signed(FMAP_9_54);
			MULT_55(8)<=signed(DIN_55_7)*signed(FMAP_9_55);
			MULT_56(8)<=signed(DIN_56_7)*signed(FMAP_9_56);
			MULT_57(8)<=signed(DIN_57_7)*signed(FMAP_9_57);
			MULT_58(8)<=signed(DIN_58_7)*signed(FMAP_9_58);
			MULT_59(8)<=signed(DIN_59_7)*signed(FMAP_9_59);
			MULT_60(8)<=signed(DIN_60_7)*signed(FMAP_9_60);
			MULT_61(8)<=signed(DIN_61_7)*signed(FMAP_9_61);
			MULT_62(8)<=signed(DIN_62_7)*signed(FMAP_9_62);
			MULT_63(8)<=signed(DIN_63_7)*signed(FMAP_9_63);
			MULT_64(8)<=signed(DIN_64_7)*signed(FMAP_9_64);
			MULT_65(8)<=signed(DIN_65_7)*signed(FMAP_9_65);
			MULT_66(8)<=signed(DIN_66_7)*signed(FMAP_9_66);
			MULT_67(8)<=signed(DIN_67_7)*signed(FMAP_9_67);
			MULT_68(8)<=signed(DIN_68_7)*signed(FMAP_9_68);
			MULT_69(8)<=signed(DIN_69_7)*signed(FMAP_9_69);
			MULT_70(8)<=signed(DIN_70_7)*signed(FMAP_9_70);
			MULT_71(8)<=signed(DIN_71_7)*signed(FMAP_9_71);
			MULT_72(8)<=signed(DIN_72_7)*signed(FMAP_9_72);
			MULT_73(8)<=signed(DIN_73_7)*signed(FMAP_9_73);
			MULT_74(8)<=signed(DIN_74_7)*signed(FMAP_9_74);
			MULT_75(8)<=signed(DIN_75_7)*signed(FMAP_9_75);
			MULT_76(8)<=signed(DIN_76_7)*signed(FMAP_9_76);
			MULT_77(8)<=signed(DIN_77_7)*signed(FMAP_9_77);
			MULT_78(8)<=signed(DIN_78_7)*signed(FMAP_9_78);
			MULT_79(8)<=signed(DIN_79_7)*signed(FMAP_9_79);
			MULT_80(8)<=signed(DIN_80_7)*signed(FMAP_9_80);
			MULT_81(8)<=signed(DIN_81_7)*signed(FMAP_9_81);
			MULT_82(8)<=signed(DIN_82_7)*signed(FMAP_9_82);
			MULT_83(8)<=signed(DIN_83_7)*signed(FMAP_9_83);
			MULT_84(8)<=signed(DIN_84_7)*signed(FMAP_9_84);
			MULT_85(8)<=signed(DIN_85_7)*signed(FMAP_9_85);
			MULT_86(8)<=signed(DIN_86_7)*signed(FMAP_9_86);
			MULT_87(8)<=signed(DIN_87_7)*signed(FMAP_9_87);
			MULT_88(8)<=signed(DIN_88_7)*signed(FMAP_9_88);
			MULT_89(8)<=signed(DIN_89_7)*signed(FMAP_9_89);
			MULT_90(8)<=signed(DIN_90_7)*signed(FMAP_9_90);
			MULT_91(8)<=signed(DIN_91_7)*signed(FMAP_9_91);
			MULT_92(8)<=signed(DIN_92_7)*signed(FMAP_9_92);
			MULT_93(8)<=signed(DIN_93_7)*signed(FMAP_9_93);
			MULT_94(8)<=signed(DIN_94_7)*signed(FMAP_9_94);
			MULT_95(8)<=signed(DIN_95_7)*signed(FMAP_9_95);
			MULT_96(8)<=signed(DIN_96_7)*signed(FMAP_9_96);
			MULT_97(8)<=signed(DIN_97_7)*signed(FMAP_9_97);
			MULT_98(8)<=signed(DIN_98_7)*signed(FMAP_9_98);
			MULT_99(8)<=signed(DIN_99_7)*signed(FMAP_9_99);
			MULT_100(8)<=signed(DIN_100_7)*signed(FMAP_9_100);
			MULT_101(8)<=signed(DIN_101_7)*signed(FMAP_9_101);
			MULT_102(8)<=signed(DIN_102_7)*signed(FMAP_9_102);
			MULT_103(8)<=signed(DIN_103_7)*signed(FMAP_9_103);
			MULT_104(8)<=signed(DIN_104_7)*signed(FMAP_9_104);
			MULT_105(8)<=signed(DIN_105_7)*signed(FMAP_9_105);
			MULT_106(8)<=signed(DIN_106_7)*signed(FMAP_9_106);
			MULT_107(8)<=signed(DIN_107_7)*signed(FMAP_9_107);
			MULT_108(8)<=signed(DIN_108_7)*signed(FMAP_9_108);
			MULT_109(8)<=signed(DIN_109_7)*signed(FMAP_9_109);
			MULT_110(8)<=signed(DIN_110_7)*signed(FMAP_9_110);
			MULT_111(8)<=signed(DIN_111_7)*signed(FMAP_9_111);
			MULT_112(8)<=signed(DIN_112_7)*signed(FMAP_9_112);
			MULT_113(8)<=signed(DIN_113_7)*signed(FMAP_9_113);
			MULT_114(8)<=signed(DIN_114_7)*signed(FMAP_9_114);
			MULT_115(8)<=signed(DIN_115_7)*signed(FMAP_9_115);
			MULT_116(8)<=signed(DIN_116_7)*signed(FMAP_9_116);
			MULT_117(8)<=signed(DIN_117_7)*signed(FMAP_9_117);
			MULT_118(8)<=signed(DIN_118_7)*signed(FMAP_9_118);
			MULT_119(8)<=signed(DIN_119_7)*signed(FMAP_9_119);
			MULT_120(8)<=signed(DIN_120_7)*signed(FMAP_9_120);

			MULT_1(9)<=signed(DIN_1_7)*signed(FMAP_10_1);
			MULT_2(9)<=signed(DIN_2_7)*signed(FMAP_10_2);
			MULT_3(9)<=signed(DIN_3_7)*signed(FMAP_10_3);
			MULT_4(9)<=signed(DIN_4_7)*signed(FMAP_10_4);
			MULT_5(9)<=signed(DIN_5_7)*signed(FMAP_10_5);
			MULT_6(9)<=signed(DIN_6_7)*signed(FMAP_10_6);
			MULT_7(9)<=signed(DIN_7_7)*signed(FMAP_10_7);
			MULT_8(9)<=signed(DIN_8_7)*signed(FMAP_10_8);
			MULT_9(9)<=signed(DIN_9_7)*signed(FMAP_10_9);
			MULT_10(9)<=signed(DIN_10_7)*signed(FMAP_10_10);
			MULT_11(9)<=signed(DIN_11_7)*signed(FMAP_10_11);
			MULT_12(9)<=signed(DIN_12_7)*signed(FMAP_10_12);
			MULT_13(9)<=signed(DIN_13_7)*signed(FMAP_10_13);
			MULT_14(9)<=signed(DIN_14_7)*signed(FMAP_10_14);
			MULT_15(9)<=signed(DIN_15_7)*signed(FMAP_10_15);
			MULT_16(9)<=signed(DIN_16_7)*signed(FMAP_10_16);
			MULT_17(9)<=signed(DIN_17_7)*signed(FMAP_10_17);
			MULT_18(9)<=signed(DIN_18_7)*signed(FMAP_10_18);
			MULT_19(9)<=signed(DIN_19_7)*signed(FMAP_10_19);
			MULT_20(9)<=signed(DIN_20_7)*signed(FMAP_10_20);
			MULT_21(9)<=signed(DIN_21_7)*signed(FMAP_10_21);
			MULT_22(9)<=signed(DIN_22_7)*signed(FMAP_10_22);
			MULT_23(9)<=signed(DIN_23_7)*signed(FMAP_10_23);
			MULT_24(9)<=signed(DIN_24_7)*signed(FMAP_10_24);
			MULT_25(9)<=signed(DIN_25_7)*signed(FMAP_10_25);
			MULT_26(9)<=signed(DIN_26_7)*signed(FMAP_10_26);
			MULT_27(9)<=signed(DIN_27_7)*signed(FMAP_10_27);
			MULT_28(9)<=signed(DIN_28_7)*signed(FMAP_10_28);
			MULT_29(9)<=signed(DIN_29_7)*signed(FMAP_10_29);
			MULT_30(9)<=signed(DIN_30_7)*signed(FMAP_10_30);
			MULT_31(9)<=signed(DIN_31_7)*signed(FMAP_10_31);
			MULT_32(9)<=signed(DIN_32_7)*signed(FMAP_10_32);
			MULT_33(9)<=signed(DIN_33_7)*signed(FMAP_10_33);
			MULT_34(9)<=signed(DIN_34_7)*signed(FMAP_10_34);
			MULT_35(9)<=signed(DIN_35_7)*signed(FMAP_10_35);
			MULT_36(9)<=signed(DIN_36_7)*signed(FMAP_10_36);
			MULT_37(9)<=signed(DIN_37_7)*signed(FMAP_10_37);
			MULT_38(9)<=signed(DIN_38_7)*signed(FMAP_10_38);
			MULT_39(9)<=signed(DIN_39_7)*signed(FMAP_10_39);
			MULT_40(9)<=signed(DIN_40_7)*signed(FMAP_10_40);
			MULT_41(9)<=signed(DIN_41_7)*signed(FMAP_10_41);
			MULT_42(9)<=signed(DIN_42_7)*signed(FMAP_10_42);
			MULT_43(9)<=signed(DIN_43_7)*signed(FMAP_10_43);
			MULT_44(9)<=signed(DIN_44_7)*signed(FMAP_10_44);
			MULT_45(9)<=signed(DIN_45_7)*signed(FMAP_10_45);
			MULT_46(9)<=signed(DIN_46_7)*signed(FMAP_10_46);
			MULT_47(9)<=signed(DIN_47_7)*signed(FMAP_10_47);
			MULT_48(9)<=signed(DIN_48_7)*signed(FMAP_10_48);
			MULT_49(9)<=signed(DIN_49_7)*signed(FMAP_10_49);
			MULT_50(9)<=signed(DIN_50_7)*signed(FMAP_10_50);
			MULT_51(9)<=signed(DIN_51_7)*signed(FMAP_10_51);
			MULT_52(9)<=signed(DIN_52_7)*signed(FMAP_10_52);
			MULT_53(9)<=signed(DIN_53_7)*signed(FMAP_10_53);
			MULT_54(9)<=signed(DIN_54_7)*signed(FMAP_10_54);
			MULT_55(9)<=signed(DIN_55_7)*signed(FMAP_10_55);
			MULT_56(9)<=signed(DIN_56_7)*signed(FMAP_10_56);
			MULT_57(9)<=signed(DIN_57_7)*signed(FMAP_10_57);
			MULT_58(9)<=signed(DIN_58_7)*signed(FMAP_10_58);
			MULT_59(9)<=signed(DIN_59_7)*signed(FMAP_10_59);
			MULT_60(9)<=signed(DIN_60_7)*signed(FMAP_10_60);
			MULT_61(9)<=signed(DIN_61_7)*signed(FMAP_10_61);
			MULT_62(9)<=signed(DIN_62_7)*signed(FMAP_10_62);
			MULT_63(9)<=signed(DIN_63_7)*signed(FMAP_10_63);
			MULT_64(9)<=signed(DIN_64_7)*signed(FMAP_10_64);
			MULT_65(9)<=signed(DIN_65_7)*signed(FMAP_10_65);
			MULT_66(9)<=signed(DIN_66_7)*signed(FMAP_10_66);
			MULT_67(9)<=signed(DIN_67_7)*signed(FMAP_10_67);
			MULT_68(9)<=signed(DIN_68_7)*signed(FMAP_10_68);
			MULT_69(9)<=signed(DIN_69_7)*signed(FMAP_10_69);
			MULT_70(9)<=signed(DIN_70_7)*signed(FMAP_10_70);
			MULT_71(9)<=signed(DIN_71_7)*signed(FMAP_10_71);
			MULT_72(9)<=signed(DIN_72_7)*signed(FMAP_10_72);
			MULT_73(9)<=signed(DIN_73_7)*signed(FMAP_10_73);
			MULT_74(9)<=signed(DIN_74_7)*signed(FMAP_10_74);
			MULT_75(9)<=signed(DIN_75_7)*signed(FMAP_10_75);
			MULT_76(9)<=signed(DIN_76_7)*signed(FMAP_10_76);
			MULT_77(9)<=signed(DIN_77_7)*signed(FMAP_10_77);
			MULT_78(9)<=signed(DIN_78_7)*signed(FMAP_10_78);
			MULT_79(9)<=signed(DIN_79_7)*signed(FMAP_10_79);
			MULT_80(9)<=signed(DIN_80_7)*signed(FMAP_10_80);
			MULT_81(9)<=signed(DIN_81_7)*signed(FMAP_10_81);
			MULT_82(9)<=signed(DIN_82_7)*signed(FMAP_10_82);
			MULT_83(9)<=signed(DIN_83_7)*signed(FMAP_10_83);
			MULT_84(9)<=signed(DIN_84_7)*signed(FMAP_10_84);
			MULT_85(9)<=signed(DIN_85_7)*signed(FMAP_10_85);
			MULT_86(9)<=signed(DIN_86_7)*signed(FMAP_10_86);
			MULT_87(9)<=signed(DIN_87_7)*signed(FMAP_10_87);
			MULT_88(9)<=signed(DIN_88_7)*signed(FMAP_10_88);
			MULT_89(9)<=signed(DIN_89_7)*signed(FMAP_10_89);
			MULT_90(9)<=signed(DIN_90_7)*signed(FMAP_10_90);
			MULT_91(9)<=signed(DIN_91_7)*signed(FMAP_10_91);
			MULT_92(9)<=signed(DIN_92_7)*signed(FMAP_10_92);
			MULT_93(9)<=signed(DIN_93_7)*signed(FMAP_10_93);
			MULT_94(9)<=signed(DIN_94_7)*signed(FMAP_10_94);
			MULT_95(9)<=signed(DIN_95_7)*signed(FMAP_10_95);
			MULT_96(9)<=signed(DIN_96_7)*signed(FMAP_10_96);
			MULT_97(9)<=signed(DIN_97_7)*signed(FMAP_10_97);
			MULT_98(9)<=signed(DIN_98_7)*signed(FMAP_10_98);
			MULT_99(9)<=signed(DIN_99_7)*signed(FMAP_10_99);
			MULT_100(9)<=signed(DIN_100_7)*signed(FMAP_10_100);
			MULT_101(9)<=signed(DIN_101_7)*signed(FMAP_10_101);
			MULT_102(9)<=signed(DIN_102_7)*signed(FMAP_10_102);
			MULT_103(9)<=signed(DIN_103_7)*signed(FMAP_10_103);
			MULT_104(9)<=signed(DIN_104_7)*signed(FMAP_10_104);
			MULT_105(9)<=signed(DIN_105_7)*signed(FMAP_10_105);
			MULT_106(9)<=signed(DIN_106_7)*signed(FMAP_10_106);
			MULT_107(9)<=signed(DIN_107_7)*signed(FMAP_10_107);
			MULT_108(9)<=signed(DIN_108_7)*signed(FMAP_10_108);
			MULT_109(9)<=signed(DIN_109_7)*signed(FMAP_10_109);
			MULT_110(9)<=signed(DIN_110_7)*signed(FMAP_10_110);
			MULT_111(9)<=signed(DIN_111_7)*signed(FMAP_10_111);
			MULT_112(9)<=signed(DIN_112_7)*signed(FMAP_10_112);
			MULT_113(9)<=signed(DIN_113_7)*signed(FMAP_10_113);
			MULT_114(9)<=signed(DIN_114_7)*signed(FMAP_10_114);
			MULT_115(9)<=signed(DIN_115_7)*signed(FMAP_10_115);
			MULT_116(9)<=signed(DIN_116_7)*signed(FMAP_10_116);
			MULT_117(9)<=signed(DIN_117_7)*signed(FMAP_10_117);
			MULT_118(9)<=signed(DIN_118_7)*signed(FMAP_10_118);
			MULT_119(9)<=signed(DIN_119_7)*signed(FMAP_10_119);
			MULT_120(9)<=signed(DIN_120_7)*signed(FMAP_10_120);


                        EN_SUM_MULT_1<='1';

      -------------------------------------------- Enable MULT START --------------------------------------------				


		if EN_SUM_MULT_1 = '1' then
			------------------------------------STAGE-1--------------------------------------
			MULTS_1_1(0)<=signed(MULT_1(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(1)<=signed(MULT_1(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(2)<=signed(MULT_1(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(3)<=signed(MULT_1(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(4)<=signed(MULT_1(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(5)<=signed(MULT_1(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(6)<=signed(MULT_1(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(7)<=signed(MULT_1(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(8)<=signed(MULT_1(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_1(9)<=signed(MULT_1(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_2(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_2(0)<=signed(MULT_3(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(1)<=signed(MULT_3(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(2)<=signed(MULT_3(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(3)<=signed(MULT_3(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(4)<=signed(MULT_3(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(5)<=signed(MULT_3(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(6)<=signed(MULT_3(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(7)<=signed(MULT_3(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(8)<=signed(MULT_3(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_2(9)<=signed(MULT_3(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_4(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_3(0)<=signed(MULT_5(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(1)<=signed(MULT_5(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(2)<=signed(MULT_5(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(3)<=signed(MULT_5(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(4)<=signed(MULT_5(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(5)<=signed(MULT_5(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(6)<=signed(MULT_5(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(7)<=signed(MULT_5(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(8)<=signed(MULT_5(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_3(9)<=signed(MULT_5(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_6(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_4(0)<=signed(MULT_7(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(1)<=signed(MULT_7(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(2)<=signed(MULT_7(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(3)<=signed(MULT_7(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(4)<=signed(MULT_7(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(5)<=signed(MULT_7(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(6)<=signed(MULT_7(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(7)<=signed(MULT_7(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(8)<=signed(MULT_7(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_4(9)<=signed(MULT_7(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_8(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_5(0)<=signed(MULT_9(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(1)<=signed(MULT_9(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(2)<=signed(MULT_9(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(3)<=signed(MULT_9(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(4)<=signed(MULT_9(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(5)<=signed(MULT_9(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(6)<=signed(MULT_9(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(7)<=signed(MULT_9(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(8)<=signed(MULT_9(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_5(9)<=signed(MULT_9(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_10(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_6(0)<=signed(MULT_11(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(1)<=signed(MULT_11(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(2)<=signed(MULT_11(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(3)<=signed(MULT_11(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(4)<=signed(MULT_11(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(5)<=signed(MULT_11(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(6)<=signed(MULT_11(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(7)<=signed(MULT_11(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(8)<=signed(MULT_11(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_6(9)<=signed(MULT_11(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_12(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_7(0)<=signed(MULT_13(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(1)<=signed(MULT_13(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(2)<=signed(MULT_13(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(3)<=signed(MULT_13(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(4)<=signed(MULT_13(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(5)<=signed(MULT_13(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(6)<=signed(MULT_13(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(7)<=signed(MULT_13(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(8)<=signed(MULT_13(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_7(9)<=signed(MULT_13(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_14(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_8(0)<=signed(MULT_15(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(1)<=signed(MULT_15(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(2)<=signed(MULT_15(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(3)<=signed(MULT_15(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(4)<=signed(MULT_15(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(5)<=signed(MULT_15(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(6)<=signed(MULT_15(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(7)<=signed(MULT_15(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(8)<=signed(MULT_15(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_8(9)<=signed(MULT_15(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_16(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_9(0)<=signed(MULT_17(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(1)<=signed(MULT_17(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(2)<=signed(MULT_17(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(3)<=signed(MULT_17(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(4)<=signed(MULT_17(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(5)<=signed(MULT_17(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(6)<=signed(MULT_17(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(7)<=signed(MULT_17(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(8)<=signed(MULT_17(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_9(9)<=signed(MULT_17(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_18(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_10(0)<=signed(MULT_19(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(1)<=signed(MULT_19(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(2)<=signed(MULT_19(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(3)<=signed(MULT_19(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(4)<=signed(MULT_19(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(5)<=signed(MULT_19(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(6)<=signed(MULT_19(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(7)<=signed(MULT_19(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(8)<=signed(MULT_19(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_10(9)<=signed(MULT_19(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_20(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_11(0)<=signed(MULT_21(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(1)<=signed(MULT_21(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(2)<=signed(MULT_21(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(3)<=signed(MULT_21(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(4)<=signed(MULT_21(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(5)<=signed(MULT_21(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(6)<=signed(MULT_21(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(7)<=signed(MULT_21(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(8)<=signed(MULT_21(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_11(9)<=signed(MULT_21(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_22(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_12(0)<=signed(MULT_23(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(1)<=signed(MULT_23(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(2)<=signed(MULT_23(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(3)<=signed(MULT_23(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(4)<=signed(MULT_23(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(5)<=signed(MULT_23(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(6)<=signed(MULT_23(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(7)<=signed(MULT_23(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(8)<=signed(MULT_23(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_12(9)<=signed(MULT_23(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_24(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_13(0)<=signed(MULT_25(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(1)<=signed(MULT_25(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(2)<=signed(MULT_25(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(3)<=signed(MULT_25(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(4)<=signed(MULT_25(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(5)<=signed(MULT_25(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(6)<=signed(MULT_25(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(7)<=signed(MULT_25(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(8)<=signed(MULT_25(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_13(9)<=signed(MULT_25(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_26(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_14(0)<=signed(MULT_27(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(1)<=signed(MULT_27(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(2)<=signed(MULT_27(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(3)<=signed(MULT_27(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(4)<=signed(MULT_27(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(5)<=signed(MULT_27(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(6)<=signed(MULT_27(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(7)<=signed(MULT_27(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(8)<=signed(MULT_27(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_14(9)<=signed(MULT_27(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_28(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_15(0)<=signed(MULT_29(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(1)<=signed(MULT_29(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(2)<=signed(MULT_29(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(3)<=signed(MULT_29(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(4)<=signed(MULT_29(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(5)<=signed(MULT_29(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(6)<=signed(MULT_29(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(7)<=signed(MULT_29(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(8)<=signed(MULT_29(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_15(9)<=signed(MULT_29(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_30(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_16(0)<=signed(MULT_31(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(1)<=signed(MULT_31(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(2)<=signed(MULT_31(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(3)<=signed(MULT_31(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(4)<=signed(MULT_31(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(5)<=signed(MULT_31(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(6)<=signed(MULT_31(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(7)<=signed(MULT_31(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(8)<=signed(MULT_31(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_16(9)<=signed(MULT_31(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_32(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_17(0)<=signed(MULT_33(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(1)<=signed(MULT_33(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(2)<=signed(MULT_33(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(3)<=signed(MULT_33(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(4)<=signed(MULT_33(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(5)<=signed(MULT_33(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(6)<=signed(MULT_33(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(7)<=signed(MULT_33(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(8)<=signed(MULT_33(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_17(9)<=signed(MULT_33(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_34(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_18(0)<=signed(MULT_35(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(1)<=signed(MULT_35(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(2)<=signed(MULT_35(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(3)<=signed(MULT_35(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(4)<=signed(MULT_35(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(5)<=signed(MULT_35(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(6)<=signed(MULT_35(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(7)<=signed(MULT_35(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(8)<=signed(MULT_35(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_18(9)<=signed(MULT_35(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_36(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_19(0)<=signed(MULT_37(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(1)<=signed(MULT_37(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(2)<=signed(MULT_37(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(3)<=signed(MULT_37(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(4)<=signed(MULT_37(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(5)<=signed(MULT_37(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(6)<=signed(MULT_37(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(7)<=signed(MULT_37(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(8)<=signed(MULT_37(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_19(9)<=signed(MULT_37(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_38(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_20(0)<=signed(MULT_39(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(1)<=signed(MULT_39(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(2)<=signed(MULT_39(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(3)<=signed(MULT_39(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(4)<=signed(MULT_39(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(5)<=signed(MULT_39(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(6)<=signed(MULT_39(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(7)<=signed(MULT_39(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(8)<=signed(MULT_39(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_20(9)<=signed(MULT_39(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_40(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_21(0)<=signed(MULT_41(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(1)<=signed(MULT_41(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(2)<=signed(MULT_41(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(3)<=signed(MULT_41(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(4)<=signed(MULT_41(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(5)<=signed(MULT_41(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(6)<=signed(MULT_41(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(7)<=signed(MULT_41(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(8)<=signed(MULT_41(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_21(9)<=signed(MULT_41(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_42(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_22(0)<=signed(MULT_43(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(1)<=signed(MULT_43(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(2)<=signed(MULT_43(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(3)<=signed(MULT_43(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(4)<=signed(MULT_43(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(5)<=signed(MULT_43(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(6)<=signed(MULT_43(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(7)<=signed(MULT_43(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(8)<=signed(MULT_43(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_22(9)<=signed(MULT_43(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_44(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_23(0)<=signed(MULT_45(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(1)<=signed(MULT_45(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(2)<=signed(MULT_45(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(3)<=signed(MULT_45(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(4)<=signed(MULT_45(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(5)<=signed(MULT_45(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(6)<=signed(MULT_45(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(7)<=signed(MULT_45(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(8)<=signed(MULT_45(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_23(9)<=signed(MULT_45(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_46(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_24(0)<=signed(MULT_47(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(1)<=signed(MULT_47(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(2)<=signed(MULT_47(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(3)<=signed(MULT_47(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(4)<=signed(MULT_47(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(5)<=signed(MULT_47(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(6)<=signed(MULT_47(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(7)<=signed(MULT_47(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(8)<=signed(MULT_47(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_24(9)<=signed(MULT_47(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_48(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_25(0)<=signed(MULT_49(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(1)<=signed(MULT_49(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(2)<=signed(MULT_49(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(3)<=signed(MULT_49(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(4)<=signed(MULT_49(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(5)<=signed(MULT_49(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(6)<=signed(MULT_49(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(7)<=signed(MULT_49(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(8)<=signed(MULT_49(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_25(9)<=signed(MULT_49(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_50(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_26(0)<=signed(MULT_51(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(1)<=signed(MULT_51(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(2)<=signed(MULT_51(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(3)<=signed(MULT_51(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(4)<=signed(MULT_51(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(5)<=signed(MULT_51(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(6)<=signed(MULT_51(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(7)<=signed(MULT_51(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(8)<=signed(MULT_51(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_26(9)<=signed(MULT_51(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_52(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_27(0)<=signed(MULT_53(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(1)<=signed(MULT_53(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(2)<=signed(MULT_53(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(3)<=signed(MULT_53(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(4)<=signed(MULT_53(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(5)<=signed(MULT_53(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(6)<=signed(MULT_53(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(7)<=signed(MULT_53(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(8)<=signed(MULT_53(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_27(9)<=signed(MULT_53(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_54(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_28(0)<=signed(MULT_55(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(1)<=signed(MULT_55(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(2)<=signed(MULT_55(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(3)<=signed(MULT_55(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(4)<=signed(MULT_55(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(5)<=signed(MULT_55(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(6)<=signed(MULT_55(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(7)<=signed(MULT_55(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(8)<=signed(MULT_55(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_28(9)<=signed(MULT_55(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_56(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_29(0)<=signed(MULT_57(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(1)<=signed(MULT_57(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(2)<=signed(MULT_57(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(3)<=signed(MULT_57(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(4)<=signed(MULT_57(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(5)<=signed(MULT_57(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(6)<=signed(MULT_57(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(7)<=signed(MULT_57(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(8)<=signed(MULT_57(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_29(9)<=signed(MULT_57(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_58(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_30(0)<=signed(MULT_59(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(1)<=signed(MULT_59(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(2)<=signed(MULT_59(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(3)<=signed(MULT_59(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(4)<=signed(MULT_59(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(5)<=signed(MULT_59(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(6)<=signed(MULT_59(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(7)<=signed(MULT_59(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(8)<=signed(MULT_59(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_30(9)<=signed(MULT_59(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_60(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_31(0)<=signed(MULT_61(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(1)<=signed(MULT_61(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(2)<=signed(MULT_61(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(3)<=signed(MULT_61(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(4)<=signed(MULT_61(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(5)<=signed(MULT_61(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(6)<=signed(MULT_61(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(7)<=signed(MULT_61(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(8)<=signed(MULT_61(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_31(9)<=signed(MULT_61(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_62(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_32(0)<=signed(MULT_63(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(1)<=signed(MULT_63(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(2)<=signed(MULT_63(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(3)<=signed(MULT_63(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(4)<=signed(MULT_63(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(5)<=signed(MULT_63(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(6)<=signed(MULT_63(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(7)<=signed(MULT_63(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(8)<=signed(MULT_63(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_32(9)<=signed(MULT_63(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_64(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_33(0)<=signed(MULT_65(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(1)<=signed(MULT_65(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(2)<=signed(MULT_65(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(3)<=signed(MULT_65(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(4)<=signed(MULT_65(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(5)<=signed(MULT_65(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(6)<=signed(MULT_65(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(7)<=signed(MULT_65(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(8)<=signed(MULT_65(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_33(9)<=signed(MULT_65(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_66(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_34(0)<=signed(MULT_67(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(1)<=signed(MULT_67(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(2)<=signed(MULT_67(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(3)<=signed(MULT_67(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(4)<=signed(MULT_67(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(5)<=signed(MULT_67(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(6)<=signed(MULT_67(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(7)<=signed(MULT_67(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(8)<=signed(MULT_67(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_34(9)<=signed(MULT_67(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_68(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_35(0)<=signed(MULT_69(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(1)<=signed(MULT_69(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(2)<=signed(MULT_69(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(3)<=signed(MULT_69(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(4)<=signed(MULT_69(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(5)<=signed(MULT_69(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(6)<=signed(MULT_69(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(7)<=signed(MULT_69(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(8)<=signed(MULT_69(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_35(9)<=signed(MULT_69(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_70(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_36(0)<=signed(MULT_71(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(1)<=signed(MULT_71(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(2)<=signed(MULT_71(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(3)<=signed(MULT_71(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(4)<=signed(MULT_71(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(5)<=signed(MULT_71(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(6)<=signed(MULT_71(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(7)<=signed(MULT_71(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(8)<=signed(MULT_71(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_36(9)<=signed(MULT_71(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_72(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_37(0)<=signed(MULT_73(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(1)<=signed(MULT_73(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(2)<=signed(MULT_73(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(3)<=signed(MULT_73(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(4)<=signed(MULT_73(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(5)<=signed(MULT_73(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(6)<=signed(MULT_73(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(7)<=signed(MULT_73(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(8)<=signed(MULT_73(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_37(9)<=signed(MULT_73(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_74(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_38(0)<=signed(MULT_75(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(1)<=signed(MULT_75(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(2)<=signed(MULT_75(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(3)<=signed(MULT_75(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(4)<=signed(MULT_75(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(5)<=signed(MULT_75(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(6)<=signed(MULT_75(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(7)<=signed(MULT_75(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(8)<=signed(MULT_75(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_38(9)<=signed(MULT_75(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_76(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_39(0)<=signed(MULT_77(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(1)<=signed(MULT_77(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(2)<=signed(MULT_77(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(3)<=signed(MULT_77(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(4)<=signed(MULT_77(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(5)<=signed(MULT_77(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(6)<=signed(MULT_77(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(7)<=signed(MULT_77(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(8)<=signed(MULT_77(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_39(9)<=signed(MULT_77(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_78(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_40(0)<=signed(MULT_79(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(1)<=signed(MULT_79(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(2)<=signed(MULT_79(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(3)<=signed(MULT_79(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(4)<=signed(MULT_79(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(5)<=signed(MULT_79(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(6)<=signed(MULT_79(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(7)<=signed(MULT_79(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(8)<=signed(MULT_79(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_40(9)<=signed(MULT_79(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_80(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_41(0)<=signed(MULT_81(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(1)<=signed(MULT_81(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(2)<=signed(MULT_81(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(3)<=signed(MULT_81(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(4)<=signed(MULT_81(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(5)<=signed(MULT_81(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(6)<=signed(MULT_81(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(7)<=signed(MULT_81(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(8)<=signed(MULT_81(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_41(9)<=signed(MULT_81(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_82(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_42(0)<=signed(MULT_83(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(1)<=signed(MULT_83(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(2)<=signed(MULT_83(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(3)<=signed(MULT_83(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(4)<=signed(MULT_83(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(5)<=signed(MULT_83(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(6)<=signed(MULT_83(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(7)<=signed(MULT_83(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(8)<=signed(MULT_83(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_42(9)<=signed(MULT_83(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_84(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_43(0)<=signed(MULT_85(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(1)<=signed(MULT_85(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(2)<=signed(MULT_85(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(3)<=signed(MULT_85(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(4)<=signed(MULT_85(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(5)<=signed(MULT_85(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(6)<=signed(MULT_85(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(7)<=signed(MULT_85(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(8)<=signed(MULT_85(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_43(9)<=signed(MULT_85(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_86(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_44(0)<=signed(MULT_87(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(1)<=signed(MULT_87(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(2)<=signed(MULT_87(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(3)<=signed(MULT_87(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(4)<=signed(MULT_87(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(5)<=signed(MULT_87(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(6)<=signed(MULT_87(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(7)<=signed(MULT_87(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(8)<=signed(MULT_87(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_44(9)<=signed(MULT_87(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_88(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_45(0)<=signed(MULT_89(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(1)<=signed(MULT_89(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(2)<=signed(MULT_89(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(3)<=signed(MULT_89(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(4)<=signed(MULT_89(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(5)<=signed(MULT_89(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(6)<=signed(MULT_89(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(7)<=signed(MULT_89(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(8)<=signed(MULT_89(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_45(9)<=signed(MULT_89(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_90(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_46(0)<=signed(MULT_91(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(1)<=signed(MULT_91(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(2)<=signed(MULT_91(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(3)<=signed(MULT_91(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(4)<=signed(MULT_91(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(5)<=signed(MULT_91(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(6)<=signed(MULT_91(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(7)<=signed(MULT_91(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(8)<=signed(MULT_91(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_46(9)<=signed(MULT_91(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_92(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_47(0)<=signed(MULT_93(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(1)<=signed(MULT_93(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(2)<=signed(MULT_93(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(3)<=signed(MULT_93(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(4)<=signed(MULT_93(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(5)<=signed(MULT_93(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(6)<=signed(MULT_93(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(7)<=signed(MULT_93(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(8)<=signed(MULT_93(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_47(9)<=signed(MULT_93(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_94(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_48(0)<=signed(MULT_95(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(1)<=signed(MULT_95(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(2)<=signed(MULT_95(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(3)<=signed(MULT_95(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(4)<=signed(MULT_95(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(5)<=signed(MULT_95(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(6)<=signed(MULT_95(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(7)<=signed(MULT_95(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(8)<=signed(MULT_95(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_48(9)<=signed(MULT_95(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_96(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_49(0)<=signed(MULT_97(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(1)<=signed(MULT_97(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(2)<=signed(MULT_97(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(3)<=signed(MULT_97(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(4)<=signed(MULT_97(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(5)<=signed(MULT_97(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(6)<=signed(MULT_97(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(7)<=signed(MULT_97(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(8)<=signed(MULT_97(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_49(9)<=signed(MULT_97(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_98(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_50(0)<=signed(MULT_99(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(1)<=signed(MULT_99(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(2)<=signed(MULT_99(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(3)<=signed(MULT_99(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(4)<=signed(MULT_99(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(5)<=signed(MULT_99(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(6)<=signed(MULT_99(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(7)<=signed(MULT_99(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(8)<=signed(MULT_99(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_50(9)<=signed(MULT_99(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_100(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_51(0)<=signed(MULT_101(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(1)<=signed(MULT_101(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(2)<=signed(MULT_101(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(3)<=signed(MULT_101(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(4)<=signed(MULT_101(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(5)<=signed(MULT_101(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(6)<=signed(MULT_101(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(7)<=signed(MULT_101(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(8)<=signed(MULT_101(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_51(9)<=signed(MULT_101(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_102(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_52(0)<=signed(MULT_103(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(1)<=signed(MULT_103(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(2)<=signed(MULT_103(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(3)<=signed(MULT_103(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(4)<=signed(MULT_103(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(5)<=signed(MULT_103(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(6)<=signed(MULT_103(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(7)<=signed(MULT_103(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(8)<=signed(MULT_103(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_52(9)<=signed(MULT_103(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_104(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_53(0)<=signed(MULT_105(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(1)<=signed(MULT_105(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(2)<=signed(MULT_105(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(3)<=signed(MULT_105(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(4)<=signed(MULT_105(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(5)<=signed(MULT_105(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(6)<=signed(MULT_105(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(7)<=signed(MULT_105(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(8)<=signed(MULT_105(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_53(9)<=signed(MULT_105(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_106(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_54(0)<=signed(MULT_107(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(1)<=signed(MULT_107(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(2)<=signed(MULT_107(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(3)<=signed(MULT_107(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(4)<=signed(MULT_107(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(5)<=signed(MULT_107(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(6)<=signed(MULT_107(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(7)<=signed(MULT_107(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(8)<=signed(MULT_107(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_54(9)<=signed(MULT_107(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_108(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_55(0)<=signed(MULT_109(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(1)<=signed(MULT_109(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(2)<=signed(MULT_109(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(3)<=signed(MULT_109(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(4)<=signed(MULT_109(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(5)<=signed(MULT_109(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(6)<=signed(MULT_109(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(7)<=signed(MULT_109(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(8)<=signed(MULT_109(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_55(9)<=signed(MULT_109(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_110(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_56(0)<=signed(MULT_111(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(1)<=signed(MULT_111(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(2)<=signed(MULT_111(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(3)<=signed(MULT_111(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(4)<=signed(MULT_111(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(5)<=signed(MULT_111(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(6)<=signed(MULT_111(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(7)<=signed(MULT_111(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(8)<=signed(MULT_111(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_56(9)<=signed(MULT_111(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_112(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_57(0)<=signed(MULT_113(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(1)<=signed(MULT_113(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(2)<=signed(MULT_113(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(3)<=signed(MULT_113(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(4)<=signed(MULT_113(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(5)<=signed(MULT_113(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(6)<=signed(MULT_113(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(7)<=signed(MULT_113(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(8)<=signed(MULT_113(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_57(9)<=signed(MULT_113(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_114(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_58(0)<=signed(MULT_115(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(1)<=signed(MULT_115(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(2)<=signed(MULT_115(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(3)<=signed(MULT_115(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(4)<=signed(MULT_115(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(5)<=signed(MULT_115(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(6)<=signed(MULT_115(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(7)<=signed(MULT_115(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(8)<=signed(MULT_115(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_58(9)<=signed(MULT_115(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_116(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_59(0)<=signed(MULT_117(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(1)<=signed(MULT_117(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(2)<=signed(MULT_117(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(3)<=signed(MULT_117(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(4)<=signed(MULT_117(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(5)<=signed(MULT_117(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(6)<=signed(MULT_117(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(7)<=signed(MULT_117(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(8)<=signed(MULT_117(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_59(9)<=signed(MULT_117(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_118(9)(MULT_SIZE-1-WHOLE downto DECIMAL));

			MULTS_1_60(0)<=signed(MULT_119(0)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(0)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(1)<=signed(MULT_119(1)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(1)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(2)<=signed(MULT_119(2)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(2)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(3)<=signed(MULT_119(3)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(3)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(4)<=signed(MULT_119(4)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(4)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(5)<=signed(MULT_119(5)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(5)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(6)<=signed(MULT_119(6)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(6)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(7)<=signed(MULT_119(7)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(7)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(8)<=signed(MULT_119(8)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(8)(MULT_SIZE-1-WHOLE downto DECIMAL));
			MULTS_1_60(9)<=signed(MULT_119(9)(MULT_SIZE-1-WHOLE downto DECIMAL))+signed(MULT_120(9)(MULT_SIZE-1-WHOLE downto DECIMAL));



                     EN_SUM_MULT_2<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_2 = '1' then
			------------------------------------STAGE-2--------------------------------------
			MULTS_2_1(0)<=signed(MULTS_1_1(0)(PRECISION-1 downto 0))+signed(MULTS_1_2(0)(PRECISION-1 downto 0));
			MULTS_2_1(1)<=signed(MULTS_1_1(1)(PRECISION-1 downto 0))+signed(MULTS_1_2(1)(PRECISION-1 downto 0));
			MULTS_2_1(2)<=signed(MULTS_1_1(2)(PRECISION-1 downto 0))+signed(MULTS_1_2(2)(PRECISION-1 downto 0));
			MULTS_2_1(3)<=signed(MULTS_1_1(3)(PRECISION-1 downto 0))+signed(MULTS_1_2(3)(PRECISION-1 downto 0));
			MULTS_2_1(4)<=signed(MULTS_1_1(4)(PRECISION-1 downto 0))+signed(MULTS_1_2(4)(PRECISION-1 downto 0));
			MULTS_2_1(5)<=signed(MULTS_1_1(5)(PRECISION-1 downto 0))+signed(MULTS_1_2(5)(PRECISION-1 downto 0));
			MULTS_2_1(6)<=signed(MULTS_1_1(6)(PRECISION-1 downto 0))+signed(MULTS_1_2(6)(PRECISION-1 downto 0));
			MULTS_2_1(7)<=signed(MULTS_1_1(7)(PRECISION-1 downto 0))+signed(MULTS_1_2(7)(PRECISION-1 downto 0));
			MULTS_2_1(8)<=signed(MULTS_1_1(8)(PRECISION-1 downto 0))+signed(MULTS_1_2(8)(PRECISION-1 downto 0));
			MULTS_2_1(9)<=signed(MULTS_1_1(9)(PRECISION-1 downto 0))+signed(MULTS_1_2(9)(PRECISION-1 downto 0));

			MULTS_2_2(0)<=signed(MULTS_1_3(0)(PRECISION-1 downto 0))+signed(MULTS_1_4(0)(PRECISION-1 downto 0));
			MULTS_2_2(1)<=signed(MULTS_1_3(1)(PRECISION-1 downto 0))+signed(MULTS_1_4(1)(PRECISION-1 downto 0));
			MULTS_2_2(2)<=signed(MULTS_1_3(2)(PRECISION-1 downto 0))+signed(MULTS_1_4(2)(PRECISION-1 downto 0));
			MULTS_2_2(3)<=signed(MULTS_1_3(3)(PRECISION-1 downto 0))+signed(MULTS_1_4(3)(PRECISION-1 downto 0));
			MULTS_2_2(4)<=signed(MULTS_1_3(4)(PRECISION-1 downto 0))+signed(MULTS_1_4(4)(PRECISION-1 downto 0));
			MULTS_2_2(5)<=signed(MULTS_1_3(5)(PRECISION-1 downto 0))+signed(MULTS_1_4(5)(PRECISION-1 downto 0));
			MULTS_2_2(6)<=signed(MULTS_1_3(6)(PRECISION-1 downto 0))+signed(MULTS_1_4(6)(PRECISION-1 downto 0));
			MULTS_2_2(7)<=signed(MULTS_1_3(7)(PRECISION-1 downto 0))+signed(MULTS_1_4(7)(PRECISION-1 downto 0));
			MULTS_2_2(8)<=signed(MULTS_1_3(8)(PRECISION-1 downto 0))+signed(MULTS_1_4(8)(PRECISION-1 downto 0));
			MULTS_2_2(9)<=signed(MULTS_1_3(9)(PRECISION-1 downto 0))+signed(MULTS_1_4(9)(PRECISION-1 downto 0));

			MULTS_2_3(0)<=signed(MULTS_1_5(0)(PRECISION-1 downto 0))+signed(MULTS_1_6(0)(PRECISION-1 downto 0));
			MULTS_2_3(1)<=signed(MULTS_1_5(1)(PRECISION-1 downto 0))+signed(MULTS_1_6(1)(PRECISION-1 downto 0));
			MULTS_2_3(2)<=signed(MULTS_1_5(2)(PRECISION-1 downto 0))+signed(MULTS_1_6(2)(PRECISION-1 downto 0));
			MULTS_2_3(3)<=signed(MULTS_1_5(3)(PRECISION-1 downto 0))+signed(MULTS_1_6(3)(PRECISION-1 downto 0));
			MULTS_2_3(4)<=signed(MULTS_1_5(4)(PRECISION-1 downto 0))+signed(MULTS_1_6(4)(PRECISION-1 downto 0));
			MULTS_2_3(5)<=signed(MULTS_1_5(5)(PRECISION-1 downto 0))+signed(MULTS_1_6(5)(PRECISION-1 downto 0));
			MULTS_2_3(6)<=signed(MULTS_1_5(6)(PRECISION-1 downto 0))+signed(MULTS_1_6(6)(PRECISION-1 downto 0));
			MULTS_2_3(7)<=signed(MULTS_1_5(7)(PRECISION-1 downto 0))+signed(MULTS_1_6(7)(PRECISION-1 downto 0));
			MULTS_2_3(8)<=signed(MULTS_1_5(8)(PRECISION-1 downto 0))+signed(MULTS_1_6(8)(PRECISION-1 downto 0));
			MULTS_2_3(9)<=signed(MULTS_1_5(9)(PRECISION-1 downto 0))+signed(MULTS_1_6(9)(PRECISION-1 downto 0));

			MULTS_2_4(0)<=signed(MULTS_1_7(0)(PRECISION-1 downto 0))+signed(MULTS_1_8(0)(PRECISION-1 downto 0));
			MULTS_2_4(1)<=signed(MULTS_1_7(1)(PRECISION-1 downto 0))+signed(MULTS_1_8(1)(PRECISION-1 downto 0));
			MULTS_2_4(2)<=signed(MULTS_1_7(2)(PRECISION-1 downto 0))+signed(MULTS_1_8(2)(PRECISION-1 downto 0));
			MULTS_2_4(3)<=signed(MULTS_1_7(3)(PRECISION-1 downto 0))+signed(MULTS_1_8(3)(PRECISION-1 downto 0));
			MULTS_2_4(4)<=signed(MULTS_1_7(4)(PRECISION-1 downto 0))+signed(MULTS_1_8(4)(PRECISION-1 downto 0));
			MULTS_2_4(5)<=signed(MULTS_1_7(5)(PRECISION-1 downto 0))+signed(MULTS_1_8(5)(PRECISION-1 downto 0));
			MULTS_2_4(6)<=signed(MULTS_1_7(6)(PRECISION-1 downto 0))+signed(MULTS_1_8(6)(PRECISION-1 downto 0));
			MULTS_2_4(7)<=signed(MULTS_1_7(7)(PRECISION-1 downto 0))+signed(MULTS_1_8(7)(PRECISION-1 downto 0));
			MULTS_2_4(8)<=signed(MULTS_1_7(8)(PRECISION-1 downto 0))+signed(MULTS_1_8(8)(PRECISION-1 downto 0));
			MULTS_2_4(9)<=signed(MULTS_1_7(9)(PRECISION-1 downto 0))+signed(MULTS_1_8(9)(PRECISION-1 downto 0));

			MULTS_2_5(0)<=signed(MULTS_1_9(0)(PRECISION-1 downto 0))+signed(MULTS_1_10(0)(PRECISION-1 downto 0));
			MULTS_2_5(1)<=signed(MULTS_1_9(1)(PRECISION-1 downto 0))+signed(MULTS_1_10(1)(PRECISION-1 downto 0));
			MULTS_2_5(2)<=signed(MULTS_1_9(2)(PRECISION-1 downto 0))+signed(MULTS_1_10(2)(PRECISION-1 downto 0));
			MULTS_2_5(3)<=signed(MULTS_1_9(3)(PRECISION-1 downto 0))+signed(MULTS_1_10(3)(PRECISION-1 downto 0));
			MULTS_2_5(4)<=signed(MULTS_1_9(4)(PRECISION-1 downto 0))+signed(MULTS_1_10(4)(PRECISION-1 downto 0));
			MULTS_2_5(5)<=signed(MULTS_1_9(5)(PRECISION-1 downto 0))+signed(MULTS_1_10(5)(PRECISION-1 downto 0));
			MULTS_2_5(6)<=signed(MULTS_1_9(6)(PRECISION-1 downto 0))+signed(MULTS_1_10(6)(PRECISION-1 downto 0));
			MULTS_2_5(7)<=signed(MULTS_1_9(7)(PRECISION-1 downto 0))+signed(MULTS_1_10(7)(PRECISION-1 downto 0));
			MULTS_2_5(8)<=signed(MULTS_1_9(8)(PRECISION-1 downto 0))+signed(MULTS_1_10(8)(PRECISION-1 downto 0));
			MULTS_2_5(9)<=signed(MULTS_1_9(9)(PRECISION-1 downto 0))+signed(MULTS_1_10(9)(PRECISION-1 downto 0));

			MULTS_2_6(0)<=signed(MULTS_1_11(0)(PRECISION-1 downto 0))+signed(MULTS_1_12(0)(PRECISION-1 downto 0));
			MULTS_2_6(1)<=signed(MULTS_1_11(1)(PRECISION-1 downto 0))+signed(MULTS_1_12(1)(PRECISION-1 downto 0));
			MULTS_2_6(2)<=signed(MULTS_1_11(2)(PRECISION-1 downto 0))+signed(MULTS_1_12(2)(PRECISION-1 downto 0));
			MULTS_2_6(3)<=signed(MULTS_1_11(3)(PRECISION-1 downto 0))+signed(MULTS_1_12(3)(PRECISION-1 downto 0));
			MULTS_2_6(4)<=signed(MULTS_1_11(4)(PRECISION-1 downto 0))+signed(MULTS_1_12(4)(PRECISION-1 downto 0));
			MULTS_2_6(5)<=signed(MULTS_1_11(5)(PRECISION-1 downto 0))+signed(MULTS_1_12(5)(PRECISION-1 downto 0));
			MULTS_2_6(6)<=signed(MULTS_1_11(6)(PRECISION-1 downto 0))+signed(MULTS_1_12(6)(PRECISION-1 downto 0));
			MULTS_2_6(7)<=signed(MULTS_1_11(7)(PRECISION-1 downto 0))+signed(MULTS_1_12(7)(PRECISION-1 downto 0));
			MULTS_2_6(8)<=signed(MULTS_1_11(8)(PRECISION-1 downto 0))+signed(MULTS_1_12(8)(PRECISION-1 downto 0));
			MULTS_2_6(9)<=signed(MULTS_1_11(9)(PRECISION-1 downto 0))+signed(MULTS_1_12(9)(PRECISION-1 downto 0));

			MULTS_2_7(0)<=signed(MULTS_1_13(0)(PRECISION-1 downto 0))+signed(MULTS_1_14(0)(PRECISION-1 downto 0));
			MULTS_2_7(1)<=signed(MULTS_1_13(1)(PRECISION-1 downto 0))+signed(MULTS_1_14(1)(PRECISION-1 downto 0));
			MULTS_2_7(2)<=signed(MULTS_1_13(2)(PRECISION-1 downto 0))+signed(MULTS_1_14(2)(PRECISION-1 downto 0));
			MULTS_2_7(3)<=signed(MULTS_1_13(3)(PRECISION-1 downto 0))+signed(MULTS_1_14(3)(PRECISION-1 downto 0));
			MULTS_2_7(4)<=signed(MULTS_1_13(4)(PRECISION-1 downto 0))+signed(MULTS_1_14(4)(PRECISION-1 downto 0));
			MULTS_2_7(5)<=signed(MULTS_1_13(5)(PRECISION-1 downto 0))+signed(MULTS_1_14(5)(PRECISION-1 downto 0));
			MULTS_2_7(6)<=signed(MULTS_1_13(6)(PRECISION-1 downto 0))+signed(MULTS_1_14(6)(PRECISION-1 downto 0));
			MULTS_2_7(7)<=signed(MULTS_1_13(7)(PRECISION-1 downto 0))+signed(MULTS_1_14(7)(PRECISION-1 downto 0));
			MULTS_2_7(8)<=signed(MULTS_1_13(8)(PRECISION-1 downto 0))+signed(MULTS_1_14(8)(PRECISION-1 downto 0));
			MULTS_2_7(9)<=signed(MULTS_1_13(9)(PRECISION-1 downto 0))+signed(MULTS_1_14(9)(PRECISION-1 downto 0));

			MULTS_2_8(0)<=signed(MULTS_1_15(0)(PRECISION-1 downto 0))+signed(MULTS_1_16(0)(PRECISION-1 downto 0));
			MULTS_2_8(1)<=signed(MULTS_1_15(1)(PRECISION-1 downto 0))+signed(MULTS_1_16(1)(PRECISION-1 downto 0));
			MULTS_2_8(2)<=signed(MULTS_1_15(2)(PRECISION-1 downto 0))+signed(MULTS_1_16(2)(PRECISION-1 downto 0));
			MULTS_2_8(3)<=signed(MULTS_1_15(3)(PRECISION-1 downto 0))+signed(MULTS_1_16(3)(PRECISION-1 downto 0));
			MULTS_2_8(4)<=signed(MULTS_1_15(4)(PRECISION-1 downto 0))+signed(MULTS_1_16(4)(PRECISION-1 downto 0));
			MULTS_2_8(5)<=signed(MULTS_1_15(5)(PRECISION-1 downto 0))+signed(MULTS_1_16(5)(PRECISION-1 downto 0));
			MULTS_2_8(6)<=signed(MULTS_1_15(6)(PRECISION-1 downto 0))+signed(MULTS_1_16(6)(PRECISION-1 downto 0));
			MULTS_2_8(7)<=signed(MULTS_1_15(7)(PRECISION-1 downto 0))+signed(MULTS_1_16(7)(PRECISION-1 downto 0));
			MULTS_2_8(8)<=signed(MULTS_1_15(8)(PRECISION-1 downto 0))+signed(MULTS_1_16(8)(PRECISION-1 downto 0));
			MULTS_2_8(9)<=signed(MULTS_1_15(9)(PRECISION-1 downto 0))+signed(MULTS_1_16(9)(PRECISION-1 downto 0));

			MULTS_2_9(0)<=signed(MULTS_1_17(0)(PRECISION-1 downto 0))+signed(MULTS_1_18(0)(PRECISION-1 downto 0));
			MULTS_2_9(1)<=signed(MULTS_1_17(1)(PRECISION-1 downto 0))+signed(MULTS_1_18(1)(PRECISION-1 downto 0));
			MULTS_2_9(2)<=signed(MULTS_1_17(2)(PRECISION-1 downto 0))+signed(MULTS_1_18(2)(PRECISION-1 downto 0));
			MULTS_2_9(3)<=signed(MULTS_1_17(3)(PRECISION-1 downto 0))+signed(MULTS_1_18(3)(PRECISION-1 downto 0));
			MULTS_2_9(4)<=signed(MULTS_1_17(4)(PRECISION-1 downto 0))+signed(MULTS_1_18(4)(PRECISION-1 downto 0));
			MULTS_2_9(5)<=signed(MULTS_1_17(5)(PRECISION-1 downto 0))+signed(MULTS_1_18(5)(PRECISION-1 downto 0));
			MULTS_2_9(6)<=signed(MULTS_1_17(6)(PRECISION-1 downto 0))+signed(MULTS_1_18(6)(PRECISION-1 downto 0));
			MULTS_2_9(7)<=signed(MULTS_1_17(7)(PRECISION-1 downto 0))+signed(MULTS_1_18(7)(PRECISION-1 downto 0));
			MULTS_2_9(8)<=signed(MULTS_1_17(8)(PRECISION-1 downto 0))+signed(MULTS_1_18(8)(PRECISION-1 downto 0));
			MULTS_2_9(9)<=signed(MULTS_1_17(9)(PRECISION-1 downto 0))+signed(MULTS_1_18(9)(PRECISION-1 downto 0));

			MULTS_2_10(0)<=signed(MULTS_1_19(0)(PRECISION-1 downto 0))+signed(MULTS_1_20(0)(PRECISION-1 downto 0));
			MULTS_2_10(1)<=signed(MULTS_1_19(1)(PRECISION-1 downto 0))+signed(MULTS_1_20(1)(PRECISION-1 downto 0));
			MULTS_2_10(2)<=signed(MULTS_1_19(2)(PRECISION-1 downto 0))+signed(MULTS_1_20(2)(PRECISION-1 downto 0));
			MULTS_2_10(3)<=signed(MULTS_1_19(3)(PRECISION-1 downto 0))+signed(MULTS_1_20(3)(PRECISION-1 downto 0));
			MULTS_2_10(4)<=signed(MULTS_1_19(4)(PRECISION-1 downto 0))+signed(MULTS_1_20(4)(PRECISION-1 downto 0));
			MULTS_2_10(5)<=signed(MULTS_1_19(5)(PRECISION-1 downto 0))+signed(MULTS_1_20(5)(PRECISION-1 downto 0));
			MULTS_2_10(6)<=signed(MULTS_1_19(6)(PRECISION-1 downto 0))+signed(MULTS_1_20(6)(PRECISION-1 downto 0));
			MULTS_2_10(7)<=signed(MULTS_1_19(7)(PRECISION-1 downto 0))+signed(MULTS_1_20(7)(PRECISION-1 downto 0));
			MULTS_2_10(8)<=signed(MULTS_1_19(8)(PRECISION-1 downto 0))+signed(MULTS_1_20(8)(PRECISION-1 downto 0));
			MULTS_2_10(9)<=signed(MULTS_1_19(9)(PRECISION-1 downto 0))+signed(MULTS_1_20(9)(PRECISION-1 downto 0));

			MULTS_2_11(0)<=signed(MULTS_1_21(0)(PRECISION-1 downto 0))+signed(MULTS_1_22(0)(PRECISION-1 downto 0));
			MULTS_2_11(1)<=signed(MULTS_1_21(1)(PRECISION-1 downto 0))+signed(MULTS_1_22(1)(PRECISION-1 downto 0));
			MULTS_2_11(2)<=signed(MULTS_1_21(2)(PRECISION-1 downto 0))+signed(MULTS_1_22(2)(PRECISION-1 downto 0));
			MULTS_2_11(3)<=signed(MULTS_1_21(3)(PRECISION-1 downto 0))+signed(MULTS_1_22(3)(PRECISION-1 downto 0));
			MULTS_2_11(4)<=signed(MULTS_1_21(4)(PRECISION-1 downto 0))+signed(MULTS_1_22(4)(PRECISION-1 downto 0));
			MULTS_2_11(5)<=signed(MULTS_1_21(5)(PRECISION-1 downto 0))+signed(MULTS_1_22(5)(PRECISION-1 downto 0));
			MULTS_2_11(6)<=signed(MULTS_1_21(6)(PRECISION-1 downto 0))+signed(MULTS_1_22(6)(PRECISION-1 downto 0));
			MULTS_2_11(7)<=signed(MULTS_1_21(7)(PRECISION-1 downto 0))+signed(MULTS_1_22(7)(PRECISION-1 downto 0));
			MULTS_2_11(8)<=signed(MULTS_1_21(8)(PRECISION-1 downto 0))+signed(MULTS_1_22(8)(PRECISION-1 downto 0));
			MULTS_2_11(9)<=signed(MULTS_1_21(9)(PRECISION-1 downto 0))+signed(MULTS_1_22(9)(PRECISION-1 downto 0));

			MULTS_2_12(0)<=signed(MULTS_1_23(0)(PRECISION-1 downto 0))+signed(MULTS_1_24(0)(PRECISION-1 downto 0));
			MULTS_2_12(1)<=signed(MULTS_1_23(1)(PRECISION-1 downto 0))+signed(MULTS_1_24(1)(PRECISION-1 downto 0));
			MULTS_2_12(2)<=signed(MULTS_1_23(2)(PRECISION-1 downto 0))+signed(MULTS_1_24(2)(PRECISION-1 downto 0));
			MULTS_2_12(3)<=signed(MULTS_1_23(3)(PRECISION-1 downto 0))+signed(MULTS_1_24(3)(PRECISION-1 downto 0));
			MULTS_2_12(4)<=signed(MULTS_1_23(4)(PRECISION-1 downto 0))+signed(MULTS_1_24(4)(PRECISION-1 downto 0));
			MULTS_2_12(5)<=signed(MULTS_1_23(5)(PRECISION-1 downto 0))+signed(MULTS_1_24(5)(PRECISION-1 downto 0));
			MULTS_2_12(6)<=signed(MULTS_1_23(6)(PRECISION-1 downto 0))+signed(MULTS_1_24(6)(PRECISION-1 downto 0));
			MULTS_2_12(7)<=signed(MULTS_1_23(7)(PRECISION-1 downto 0))+signed(MULTS_1_24(7)(PRECISION-1 downto 0));
			MULTS_2_12(8)<=signed(MULTS_1_23(8)(PRECISION-1 downto 0))+signed(MULTS_1_24(8)(PRECISION-1 downto 0));
			MULTS_2_12(9)<=signed(MULTS_1_23(9)(PRECISION-1 downto 0))+signed(MULTS_1_24(9)(PRECISION-1 downto 0));

			MULTS_2_13(0)<=signed(MULTS_1_25(0)(PRECISION-1 downto 0))+signed(MULTS_1_26(0)(PRECISION-1 downto 0));
			MULTS_2_13(1)<=signed(MULTS_1_25(1)(PRECISION-1 downto 0))+signed(MULTS_1_26(1)(PRECISION-1 downto 0));
			MULTS_2_13(2)<=signed(MULTS_1_25(2)(PRECISION-1 downto 0))+signed(MULTS_1_26(2)(PRECISION-1 downto 0));
			MULTS_2_13(3)<=signed(MULTS_1_25(3)(PRECISION-1 downto 0))+signed(MULTS_1_26(3)(PRECISION-1 downto 0));
			MULTS_2_13(4)<=signed(MULTS_1_25(4)(PRECISION-1 downto 0))+signed(MULTS_1_26(4)(PRECISION-1 downto 0));
			MULTS_2_13(5)<=signed(MULTS_1_25(5)(PRECISION-1 downto 0))+signed(MULTS_1_26(5)(PRECISION-1 downto 0));
			MULTS_2_13(6)<=signed(MULTS_1_25(6)(PRECISION-1 downto 0))+signed(MULTS_1_26(6)(PRECISION-1 downto 0));
			MULTS_2_13(7)<=signed(MULTS_1_25(7)(PRECISION-1 downto 0))+signed(MULTS_1_26(7)(PRECISION-1 downto 0));
			MULTS_2_13(8)<=signed(MULTS_1_25(8)(PRECISION-1 downto 0))+signed(MULTS_1_26(8)(PRECISION-1 downto 0));
			MULTS_2_13(9)<=signed(MULTS_1_25(9)(PRECISION-1 downto 0))+signed(MULTS_1_26(9)(PRECISION-1 downto 0));

			MULTS_2_14(0)<=signed(MULTS_1_27(0)(PRECISION-1 downto 0))+signed(MULTS_1_28(0)(PRECISION-1 downto 0));
			MULTS_2_14(1)<=signed(MULTS_1_27(1)(PRECISION-1 downto 0))+signed(MULTS_1_28(1)(PRECISION-1 downto 0));
			MULTS_2_14(2)<=signed(MULTS_1_27(2)(PRECISION-1 downto 0))+signed(MULTS_1_28(2)(PRECISION-1 downto 0));
			MULTS_2_14(3)<=signed(MULTS_1_27(3)(PRECISION-1 downto 0))+signed(MULTS_1_28(3)(PRECISION-1 downto 0));
			MULTS_2_14(4)<=signed(MULTS_1_27(4)(PRECISION-1 downto 0))+signed(MULTS_1_28(4)(PRECISION-1 downto 0));
			MULTS_2_14(5)<=signed(MULTS_1_27(5)(PRECISION-1 downto 0))+signed(MULTS_1_28(5)(PRECISION-1 downto 0));
			MULTS_2_14(6)<=signed(MULTS_1_27(6)(PRECISION-1 downto 0))+signed(MULTS_1_28(6)(PRECISION-1 downto 0));
			MULTS_2_14(7)<=signed(MULTS_1_27(7)(PRECISION-1 downto 0))+signed(MULTS_1_28(7)(PRECISION-1 downto 0));
			MULTS_2_14(8)<=signed(MULTS_1_27(8)(PRECISION-1 downto 0))+signed(MULTS_1_28(8)(PRECISION-1 downto 0));
			MULTS_2_14(9)<=signed(MULTS_1_27(9)(PRECISION-1 downto 0))+signed(MULTS_1_28(9)(PRECISION-1 downto 0));

			MULTS_2_15(0)<=signed(MULTS_1_29(0)(PRECISION-1 downto 0))+signed(MULTS_1_30(0)(PRECISION-1 downto 0));
			MULTS_2_15(1)<=signed(MULTS_1_29(1)(PRECISION-1 downto 0))+signed(MULTS_1_30(1)(PRECISION-1 downto 0));
			MULTS_2_15(2)<=signed(MULTS_1_29(2)(PRECISION-1 downto 0))+signed(MULTS_1_30(2)(PRECISION-1 downto 0));
			MULTS_2_15(3)<=signed(MULTS_1_29(3)(PRECISION-1 downto 0))+signed(MULTS_1_30(3)(PRECISION-1 downto 0));
			MULTS_2_15(4)<=signed(MULTS_1_29(4)(PRECISION-1 downto 0))+signed(MULTS_1_30(4)(PRECISION-1 downto 0));
			MULTS_2_15(5)<=signed(MULTS_1_29(5)(PRECISION-1 downto 0))+signed(MULTS_1_30(5)(PRECISION-1 downto 0));
			MULTS_2_15(6)<=signed(MULTS_1_29(6)(PRECISION-1 downto 0))+signed(MULTS_1_30(6)(PRECISION-1 downto 0));
			MULTS_2_15(7)<=signed(MULTS_1_29(7)(PRECISION-1 downto 0))+signed(MULTS_1_30(7)(PRECISION-1 downto 0));
			MULTS_2_15(8)<=signed(MULTS_1_29(8)(PRECISION-1 downto 0))+signed(MULTS_1_30(8)(PRECISION-1 downto 0));
			MULTS_2_15(9)<=signed(MULTS_1_29(9)(PRECISION-1 downto 0))+signed(MULTS_1_30(9)(PRECISION-1 downto 0));



                         EN_SUM_MULT_3<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_3 = '1' then
			------------------------------------STAGE-3--------------------------------------
			MULTS_3_1(0)<=signed(MULTS_2_1(0)(PRECISION-1 downto 0))+signed(MULTS_2_2(0)(PRECISION-1 downto 0));
			MULTS_3_1(1)<=signed(MULTS_2_1(1)(PRECISION-1 downto 0))+signed(MULTS_2_2(1)(PRECISION-1 downto 0));
			MULTS_3_1(2)<=signed(MULTS_2_1(2)(PRECISION-1 downto 0))+signed(MULTS_2_2(2)(PRECISION-1 downto 0));
			MULTS_3_1(3)<=signed(MULTS_2_1(3)(PRECISION-1 downto 0))+signed(MULTS_2_2(3)(PRECISION-1 downto 0));
			MULTS_3_1(4)<=signed(MULTS_2_1(4)(PRECISION-1 downto 0))+signed(MULTS_2_2(4)(PRECISION-1 downto 0));
			MULTS_3_1(5)<=signed(MULTS_2_1(5)(PRECISION-1 downto 0))+signed(MULTS_2_2(5)(PRECISION-1 downto 0));
			MULTS_3_1(6)<=signed(MULTS_2_1(6)(PRECISION-1 downto 0))+signed(MULTS_2_2(6)(PRECISION-1 downto 0));
			MULTS_3_1(7)<=signed(MULTS_2_1(7)(PRECISION-1 downto 0))+signed(MULTS_2_2(7)(PRECISION-1 downto 0));
			MULTS_3_1(8)<=signed(MULTS_2_1(8)(PRECISION-1 downto 0))+signed(MULTS_2_2(8)(PRECISION-1 downto 0));
			MULTS_3_1(9)<=signed(MULTS_2_1(9)(PRECISION-1 downto 0))+signed(MULTS_2_2(9)(PRECISION-1 downto 0));

			MULTS_3_2(0)<=signed(MULTS_2_3(0)(PRECISION-1 downto 0))+signed(MULTS_2_4(0)(PRECISION-1 downto 0));
			MULTS_3_2(1)<=signed(MULTS_2_3(1)(PRECISION-1 downto 0))+signed(MULTS_2_4(1)(PRECISION-1 downto 0));
			MULTS_3_2(2)<=signed(MULTS_2_3(2)(PRECISION-1 downto 0))+signed(MULTS_2_4(2)(PRECISION-1 downto 0));
			MULTS_3_2(3)<=signed(MULTS_2_3(3)(PRECISION-1 downto 0))+signed(MULTS_2_4(3)(PRECISION-1 downto 0));
			MULTS_3_2(4)<=signed(MULTS_2_3(4)(PRECISION-1 downto 0))+signed(MULTS_2_4(4)(PRECISION-1 downto 0));
			MULTS_3_2(5)<=signed(MULTS_2_3(5)(PRECISION-1 downto 0))+signed(MULTS_2_4(5)(PRECISION-1 downto 0));
			MULTS_3_2(6)<=signed(MULTS_2_3(6)(PRECISION-1 downto 0))+signed(MULTS_2_4(6)(PRECISION-1 downto 0));
			MULTS_3_2(7)<=signed(MULTS_2_3(7)(PRECISION-1 downto 0))+signed(MULTS_2_4(7)(PRECISION-1 downto 0));
			MULTS_3_2(8)<=signed(MULTS_2_3(8)(PRECISION-1 downto 0))+signed(MULTS_2_4(8)(PRECISION-1 downto 0));
			MULTS_3_2(9)<=signed(MULTS_2_3(9)(PRECISION-1 downto 0))+signed(MULTS_2_4(9)(PRECISION-1 downto 0));

			MULTS_3_3(0)<=signed(MULTS_2_5(0)(PRECISION-1 downto 0))+signed(MULTS_2_6(0)(PRECISION-1 downto 0));
			MULTS_3_3(1)<=signed(MULTS_2_5(1)(PRECISION-1 downto 0))+signed(MULTS_2_6(1)(PRECISION-1 downto 0));
			MULTS_3_3(2)<=signed(MULTS_2_5(2)(PRECISION-1 downto 0))+signed(MULTS_2_6(2)(PRECISION-1 downto 0));
			MULTS_3_3(3)<=signed(MULTS_2_5(3)(PRECISION-1 downto 0))+signed(MULTS_2_6(3)(PRECISION-1 downto 0));
			MULTS_3_3(4)<=signed(MULTS_2_5(4)(PRECISION-1 downto 0))+signed(MULTS_2_6(4)(PRECISION-1 downto 0));
			MULTS_3_3(5)<=signed(MULTS_2_5(5)(PRECISION-1 downto 0))+signed(MULTS_2_6(5)(PRECISION-1 downto 0));
			MULTS_3_3(6)<=signed(MULTS_2_5(6)(PRECISION-1 downto 0))+signed(MULTS_2_6(6)(PRECISION-1 downto 0));
			MULTS_3_3(7)<=signed(MULTS_2_5(7)(PRECISION-1 downto 0))+signed(MULTS_2_6(7)(PRECISION-1 downto 0));
			MULTS_3_3(8)<=signed(MULTS_2_5(8)(PRECISION-1 downto 0))+signed(MULTS_2_6(8)(PRECISION-1 downto 0));
			MULTS_3_3(9)<=signed(MULTS_2_5(9)(PRECISION-1 downto 0))+signed(MULTS_2_6(9)(PRECISION-1 downto 0));

			MULTS_3_4(0)<=signed(MULTS_2_7(0)(PRECISION-1 downto 0))+signed(MULTS_2_8(0)(PRECISION-1 downto 0));
			MULTS_3_4(1)<=signed(MULTS_2_7(1)(PRECISION-1 downto 0))+signed(MULTS_2_8(1)(PRECISION-1 downto 0));
			MULTS_3_4(2)<=signed(MULTS_2_7(2)(PRECISION-1 downto 0))+signed(MULTS_2_8(2)(PRECISION-1 downto 0));
			MULTS_3_4(3)<=signed(MULTS_2_7(3)(PRECISION-1 downto 0))+signed(MULTS_2_8(3)(PRECISION-1 downto 0));
			MULTS_3_4(4)<=signed(MULTS_2_7(4)(PRECISION-1 downto 0))+signed(MULTS_2_8(4)(PRECISION-1 downto 0));
			MULTS_3_4(5)<=signed(MULTS_2_7(5)(PRECISION-1 downto 0))+signed(MULTS_2_8(5)(PRECISION-1 downto 0));
			MULTS_3_4(6)<=signed(MULTS_2_7(6)(PRECISION-1 downto 0))+signed(MULTS_2_8(6)(PRECISION-1 downto 0));
			MULTS_3_4(7)<=signed(MULTS_2_7(7)(PRECISION-1 downto 0))+signed(MULTS_2_8(7)(PRECISION-1 downto 0));
			MULTS_3_4(8)<=signed(MULTS_2_7(8)(PRECISION-1 downto 0))+signed(MULTS_2_8(8)(PRECISION-1 downto 0));
			MULTS_3_4(9)<=signed(MULTS_2_7(9)(PRECISION-1 downto 0))+signed(MULTS_2_8(9)(PRECISION-1 downto 0));

			MULTS_3_5(0)<=signed(MULTS_2_9(0)(PRECISION-1 downto 0))+signed(MULTS_2_10(0)(PRECISION-1 downto 0));
			MULTS_3_5(1)<=signed(MULTS_2_9(1)(PRECISION-1 downto 0))+signed(MULTS_2_10(1)(PRECISION-1 downto 0));
			MULTS_3_5(2)<=signed(MULTS_2_9(2)(PRECISION-1 downto 0))+signed(MULTS_2_10(2)(PRECISION-1 downto 0));
			MULTS_3_5(3)<=signed(MULTS_2_9(3)(PRECISION-1 downto 0))+signed(MULTS_2_10(3)(PRECISION-1 downto 0));
			MULTS_3_5(4)<=signed(MULTS_2_9(4)(PRECISION-1 downto 0))+signed(MULTS_2_10(4)(PRECISION-1 downto 0));
			MULTS_3_5(5)<=signed(MULTS_2_9(5)(PRECISION-1 downto 0))+signed(MULTS_2_10(5)(PRECISION-1 downto 0));
			MULTS_3_5(6)<=signed(MULTS_2_9(6)(PRECISION-1 downto 0))+signed(MULTS_2_10(6)(PRECISION-1 downto 0));
			MULTS_3_5(7)<=signed(MULTS_2_9(7)(PRECISION-1 downto 0))+signed(MULTS_2_10(7)(PRECISION-1 downto 0));
			MULTS_3_5(8)<=signed(MULTS_2_9(8)(PRECISION-1 downto 0))+signed(MULTS_2_10(8)(PRECISION-1 downto 0));
			MULTS_3_5(9)<=signed(MULTS_2_9(9)(PRECISION-1 downto 0))+signed(MULTS_2_10(9)(PRECISION-1 downto 0));

			MULTS_3_6(0)<=signed(MULTS_2_11(0)(PRECISION-1 downto 0))+signed(MULTS_2_12(0)(PRECISION-1 downto 0));
			MULTS_3_6(1)<=signed(MULTS_2_11(1)(PRECISION-1 downto 0))+signed(MULTS_2_12(1)(PRECISION-1 downto 0));
			MULTS_3_6(2)<=signed(MULTS_2_11(2)(PRECISION-1 downto 0))+signed(MULTS_2_12(2)(PRECISION-1 downto 0));
			MULTS_3_6(3)<=signed(MULTS_2_11(3)(PRECISION-1 downto 0))+signed(MULTS_2_12(3)(PRECISION-1 downto 0));
			MULTS_3_6(4)<=signed(MULTS_2_11(4)(PRECISION-1 downto 0))+signed(MULTS_2_12(4)(PRECISION-1 downto 0));
			MULTS_3_6(5)<=signed(MULTS_2_11(5)(PRECISION-1 downto 0))+signed(MULTS_2_12(5)(PRECISION-1 downto 0));
			MULTS_3_6(6)<=signed(MULTS_2_11(6)(PRECISION-1 downto 0))+signed(MULTS_2_12(6)(PRECISION-1 downto 0));
			MULTS_3_6(7)<=signed(MULTS_2_11(7)(PRECISION-1 downto 0))+signed(MULTS_2_12(7)(PRECISION-1 downto 0));
			MULTS_3_6(8)<=signed(MULTS_2_11(8)(PRECISION-1 downto 0))+signed(MULTS_2_12(8)(PRECISION-1 downto 0));
			MULTS_3_6(9)<=signed(MULTS_2_11(9)(PRECISION-1 downto 0))+signed(MULTS_2_12(9)(PRECISION-1 downto 0));

			MULTS_3_7(0)<=signed(MULTS_2_13(0)(PRECISION-1 downto 0))+signed(MULTS_2_14(0)(PRECISION-1 downto 0));
			MULTS_3_7(1)<=signed(MULTS_2_13(1)(PRECISION-1 downto 0))+signed(MULTS_2_14(1)(PRECISION-1 downto 0));
			MULTS_3_7(2)<=signed(MULTS_2_13(2)(PRECISION-1 downto 0))+signed(MULTS_2_14(2)(PRECISION-1 downto 0));
			MULTS_3_7(3)<=signed(MULTS_2_13(3)(PRECISION-1 downto 0))+signed(MULTS_2_14(3)(PRECISION-1 downto 0));
			MULTS_3_7(4)<=signed(MULTS_2_13(4)(PRECISION-1 downto 0))+signed(MULTS_2_14(4)(PRECISION-1 downto 0));
			MULTS_3_7(5)<=signed(MULTS_2_13(5)(PRECISION-1 downto 0))+signed(MULTS_2_14(5)(PRECISION-1 downto 0));
			MULTS_3_7(6)<=signed(MULTS_2_13(6)(PRECISION-1 downto 0))+signed(MULTS_2_14(6)(PRECISION-1 downto 0));
			MULTS_3_7(7)<=signed(MULTS_2_13(7)(PRECISION-1 downto 0))+signed(MULTS_2_14(7)(PRECISION-1 downto 0));
			MULTS_3_7(8)<=signed(MULTS_2_13(8)(PRECISION-1 downto 0))+signed(MULTS_2_14(8)(PRECISION-1 downto 0));
			MULTS_3_7(9)<=signed(MULTS_2_13(9)(PRECISION-1 downto 0))+signed(MULTS_2_14(9)(PRECISION-1 downto 0));

			MULTS_3_8(0)<=signed(MULTS_2_15(0)(PRECISION-1 downto 0))+signed(MULTS_2_16(0)(PRECISION-1 downto 0));
			MULTS_3_8(1)<=signed(MULTS_2_15(1)(PRECISION-1 downto 0))+signed(MULTS_2_16(1)(PRECISION-1 downto 0));
			MULTS_3_8(2)<=signed(MULTS_2_15(2)(PRECISION-1 downto 0))+signed(MULTS_2_16(2)(PRECISION-1 downto 0));
			MULTS_3_8(3)<=signed(MULTS_2_15(3)(PRECISION-1 downto 0))+signed(MULTS_2_16(3)(PRECISION-1 downto 0));
			MULTS_3_8(4)<=signed(MULTS_2_15(4)(PRECISION-1 downto 0))+signed(MULTS_2_16(4)(PRECISION-1 downto 0));
			MULTS_3_8(5)<=signed(MULTS_2_15(5)(PRECISION-1 downto 0))+signed(MULTS_2_16(5)(PRECISION-1 downto 0));
			MULTS_3_8(6)<=signed(MULTS_2_15(6)(PRECISION-1 downto 0))+signed(MULTS_2_16(6)(PRECISION-1 downto 0));
			MULTS_3_8(7)<=signed(MULTS_2_15(7)(PRECISION-1 downto 0))+signed(MULTS_2_16(7)(PRECISION-1 downto 0));
			MULTS_3_8(8)<=signed(MULTS_2_15(8)(PRECISION-1 downto 0))+signed(MULTS_2_16(8)(PRECISION-1 downto 0));
			MULTS_3_8(9)<=signed(MULTS_2_15(9)(PRECISION-1 downto 0))+signed(MULTS_2_16(9)(PRECISION-1 downto 0));



                         EN_SUM_MULT_4<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_4 = '1' then
			------------------------------------STAGE-4--------------------------------------
			MULTS_4_1(0)<=signed(MULTS_3_1(0));
			MULTS_4_1(1)<=signed(MULTS_3_1(1));
			MULTS_4_1(2)<=signed(MULTS_3_1(2));
			MULTS_4_1(3)<=signed(MULTS_3_1(3));
			MULTS_4_1(4)<=signed(MULTS_3_1(4));
			MULTS_4_1(5)<=signed(MULTS_3_1(5));
			MULTS_4_1(6)<=signed(MULTS_3_1(6));
			MULTS_4_1(7)<=signed(MULTS_3_1(7));
			MULTS_4_1(8)<=signed(MULTS_3_1(8));
			MULTS_4_1(9)<=signed(MULTS_3_1(9));

			MULTS_4_2(0)<=signed(MULTS_3_2(0)(PRECISION-1 downto 0))+signed(MULTS_3_3(0)(PRECISION-1 downto 0));
			MULTS_4_2(1)<=signed(MULTS_3_2(1)(PRECISION-1 downto 0))+signed(MULTS_3_3(1)(PRECISION-1 downto 0));
			MULTS_4_2(2)<=signed(MULTS_3_2(2)(PRECISION-1 downto 0))+signed(MULTS_3_3(2)(PRECISION-1 downto 0));
			MULTS_4_2(3)<=signed(MULTS_3_2(3)(PRECISION-1 downto 0))+signed(MULTS_3_3(3)(PRECISION-1 downto 0));
			MULTS_4_2(4)<=signed(MULTS_3_2(4)(PRECISION-1 downto 0))+signed(MULTS_3_3(4)(PRECISION-1 downto 0));
			MULTS_4_2(5)<=signed(MULTS_3_2(5)(PRECISION-1 downto 0))+signed(MULTS_3_3(5)(PRECISION-1 downto 0));
			MULTS_4_2(6)<=signed(MULTS_3_2(6)(PRECISION-1 downto 0))+signed(MULTS_3_3(6)(PRECISION-1 downto 0));
			MULTS_4_2(7)<=signed(MULTS_3_2(7)(PRECISION-1 downto 0))+signed(MULTS_3_3(7)(PRECISION-1 downto 0));
			MULTS_4_2(8)<=signed(MULTS_3_2(8)(PRECISION-1 downto 0))+signed(MULTS_3_3(8)(PRECISION-1 downto 0));
			MULTS_4_2(9)<=signed(MULTS_3_2(9)(PRECISION-1 downto 0))+signed(MULTS_3_3(9)(PRECISION-1 downto 0));

			MULTS_4_3(0)<=signed(MULTS_3_4(0)(PRECISION-1 downto 0))+signed(MULTS_3_5(0)(PRECISION-1 downto 0));
			MULTS_4_3(1)<=signed(MULTS_3_4(1)(PRECISION-1 downto 0))+signed(MULTS_3_5(1)(PRECISION-1 downto 0));
			MULTS_4_3(2)<=signed(MULTS_3_4(2)(PRECISION-1 downto 0))+signed(MULTS_3_5(2)(PRECISION-1 downto 0));
			MULTS_4_3(3)<=signed(MULTS_3_4(3)(PRECISION-1 downto 0))+signed(MULTS_3_5(3)(PRECISION-1 downto 0));
			MULTS_4_3(4)<=signed(MULTS_3_4(4)(PRECISION-1 downto 0))+signed(MULTS_3_5(4)(PRECISION-1 downto 0));
			MULTS_4_3(5)<=signed(MULTS_3_4(5)(PRECISION-1 downto 0))+signed(MULTS_3_5(5)(PRECISION-1 downto 0));
			MULTS_4_3(6)<=signed(MULTS_3_4(6)(PRECISION-1 downto 0))+signed(MULTS_3_5(6)(PRECISION-1 downto 0));
			MULTS_4_3(7)<=signed(MULTS_3_4(7)(PRECISION-1 downto 0))+signed(MULTS_3_5(7)(PRECISION-1 downto 0));
			MULTS_4_3(8)<=signed(MULTS_3_4(8)(PRECISION-1 downto 0))+signed(MULTS_3_5(8)(PRECISION-1 downto 0));
			MULTS_4_3(9)<=signed(MULTS_3_4(9)(PRECISION-1 downto 0))+signed(MULTS_3_5(9)(PRECISION-1 downto 0));

			MULTS_4_4(0)<=signed(MULTS_3_6(0)(PRECISION-1 downto 0))+signed(MULTS_3_7(0)(PRECISION-1 downto 0));
			MULTS_4_4(1)<=signed(MULTS_3_6(1)(PRECISION-1 downto 0))+signed(MULTS_3_7(1)(PRECISION-1 downto 0));
			MULTS_4_4(2)<=signed(MULTS_3_6(2)(PRECISION-1 downto 0))+signed(MULTS_3_7(2)(PRECISION-1 downto 0));
			MULTS_4_4(3)<=signed(MULTS_3_6(3)(PRECISION-1 downto 0))+signed(MULTS_3_7(3)(PRECISION-1 downto 0));
			MULTS_4_4(4)<=signed(MULTS_3_6(4)(PRECISION-1 downto 0))+signed(MULTS_3_7(4)(PRECISION-1 downto 0));
			MULTS_4_4(5)<=signed(MULTS_3_6(5)(PRECISION-1 downto 0))+signed(MULTS_3_7(5)(PRECISION-1 downto 0));
			MULTS_4_4(6)<=signed(MULTS_3_6(6)(PRECISION-1 downto 0))+signed(MULTS_3_7(6)(PRECISION-1 downto 0));
			MULTS_4_4(7)<=signed(MULTS_3_6(7)(PRECISION-1 downto 0))+signed(MULTS_3_7(7)(PRECISION-1 downto 0));
			MULTS_4_4(8)<=signed(MULTS_3_6(8)(PRECISION-1 downto 0))+signed(MULTS_3_7(8)(PRECISION-1 downto 0));
			MULTS_4_4(9)<=signed(MULTS_3_6(9)(PRECISION-1 downto 0))+signed(MULTS_3_7(9)(PRECISION-1 downto 0));

			MULTS_4_5(0)<=signed(MULTS_3_8(0)(PRECISION-1 downto 0))+signed(MULTS_3_9(0)(PRECISION-1 downto 0));
			MULTS_4_5(1)<=signed(MULTS_3_8(1)(PRECISION-1 downto 0))+signed(MULTS_3_9(1)(PRECISION-1 downto 0));
			MULTS_4_5(2)<=signed(MULTS_3_8(2)(PRECISION-1 downto 0))+signed(MULTS_3_9(2)(PRECISION-1 downto 0));
			MULTS_4_5(3)<=signed(MULTS_3_8(3)(PRECISION-1 downto 0))+signed(MULTS_3_9(3)(PRECISION-1 downto 0));
			MULTS_4_5(4)<=signed(MULTS_3_8(4)(PRECISION-1 downto 0))+signed(MULTS_3_9(4)(PRECISION-1 downto 0));
			MULTS_4_5(5)<=signed(MULTS_3_8(5)(PRECISION-1 downto 0))+signed(MULTS_3_9(5)(PRECISION-1 downto 0));
			MULTS_4_5(6)<=signed(MULTS_3_8(6)(PRECISION-1 downto 0))+signed(MULTS_3_9(6)(PRECISION-1 downto 0));
			MULTS_4_5(7)<=signed(MULTS_3_8(7)(PRECISION-1 downto 0))+signed(MULTS_3_9(7)(PRECISION-1 downto 0));
			MULTS_4_5(8)<=signed(MULTS_3_8(8)(PRECISION-1 downto 0))+signed(MULTS_3_9(8)(PRECISION-1 downto 0));
			MULTS_4_5(9)<=signed(MULTS_3_8(9)(PRECISION-1 downto 0))+signed(MULTS_3_9(9)(PRECISION-1 downto 0));



                         EN_SUM_MULT_5<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_5 = '1' then
			------------------------------------STAGE-5--------------------------------------
			MULTS_5_1(0)<=signed(MULTS_4_1(0)(PRECISION-1 downto 0))+signed(MULTS_4_2(0)(PRECISION-1 downto 0));
			MULTS_5_1(1)<=signed(MULTS_4_1(1)(PRECISION-1 downto 0))+signed(MULTS_4_2(1)(PRECISION-1 downto 0));
			MULTS_5_1(2)<=signed(MULTS_4_1(2)(PRECISION-1 downto 0))+signed(MULTS_4_2(2)(PRECISION-1 downto 0));
			MULTS_5_1(3)<=signed(MULTS_4_1(3)(PRECISION-1 downto 0))+signed(MULTS_4_2(3)(PRECISION-1 downto 0));
			MULTS_5_1(4)<=signed(MULTS_4_1(4)(PRECISION-1 downto 0))+signed(MULTS_4_2(4)(PRECISION-1 downto 0));
			MULTS_5_1(5)<=signed(MULTS_4_1(5)(PRECISION-1 downto 0))+signed(MULTS_4_2(5)(PRECISION-1 downto 0));
			MULTS_5_1(6)<=signed(MULTS_4_1(6)(PRECISION-1 downto 0))+signed(MULTS_4_2(6)(PRECISION-1 downto 0));
			MULTS_5_1(7)<=signed(MULTS_4_1(7)(PRECISION-1 downto 0))+signed(MULTS_4_2(7)(PRECISION-1 downto 0));
			MULTS_5_1(8)<=signed(MULTS_4_1(8)(PRECISION-1 downto 0))+signed(MULTS_4_2(8)(PRECISION-1 downto 0));
			MULTS_5_1(9)<=signed(MULTS_4_1(9)(PRECISION-1 downto 0))+signed(MULTS_4_2(9)(PRECISION-1 downto 0));

			MULTS_5_2(0)<=signed(MULTS_4_3(0)(PRECISION-1 downto 0))+signed(MULTS_4_4(0)(PRECISION-1 downto 0));
			MULTS_5_2(1)<=signed(MULTS_4_3(1)(PRECISION-1 downto 0))+signed(MULTS_4_4(1)(PRECISION-1 downto 0));
			MULTS_5_2(2)<=signed(MULTS_4_3(2)(PRECISION-1 downto 0))+signed(MULTS_4_4(2)(PRECISION-1 downto 0));
			MULTS_5_2(3)<=signed(MULTS_4_3(3)(PRECISION-1 downto 0))+signed(MULTS_4_4(3)(PRECISION-1 downto 0));
			MULTS_5_2(4)<=signed(MULTS_4_3(4)(PRECISION-1 downto 0))+signed(MULTS_4_4(4)(PRECISION-1 downto 0));
			MULTS_5_2(5)<=signed(MULTS_4_3(5)(PRECISION-1 downto 0))+signed(MULTS_4_4(5)(PRECISION-1 downto 0));
			MULTS_5_2(6)<=signed(MULTS_4_3(6)(PRECISION-1 downto 0))+signed(MULTS_4_4(6)(PRECISION-1 downto 0));
			MULTS_5_2(7)<=signed(MULTS_4_3(7)(PRECISION-1 downto 0))+signed(MULTS_4_4(7)(PRECISION-1 downto 0));
			MULTS_5_2(8)<=signed(MULTS_4_3(8)(PRECISION-1 downto 0))+signed(MULTS_4_4(8)(PRECISION-1 downto 0));
			MULTS_5_2(9)<=signed(MULTS_4_3(9)(PRECISION-1 downto 0))+signed(MULTS_4_4(9)(PRECISION-1 downto 0));



                         EN_SUM_MULT_6<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_6 = '1' then
			------------------------------------STAGE-6--------------------------------------
			MULTS_6_1(0)<=signed(MULTS_5_1(0)(PRECISION-1 downto 0))+signed(MULTS_5_2(0)(PRECISION-1 downto 0));
			MULTS_6_1(1)<=signed(MULTS_5_1(1)(PRECISION-1 downto 0))+signed(MULTS_5_2(1)(PRECISION-1 downto 0));
			MULTS_6_1(2)<=signed(MULTS_5_1(2)(PRECISION-1 downto 0))+signed(MULTS_5_2(2)(PRECISION-1 downto 0));
			MULTS_6_1(3)<=signed(MULTS_5_1(3)(PRECISION-1 downto 0))+signed(MULTS_5_2(3)(PRECISION-1 downto 0));
			MULTS_6_1(4)<=signed(MULTS_5_1(4)(PRECISION-1 downto 0))+signed(MULTS_5_2(4)(PRECISION-1 downto 0));
			MULTS_6_1(5)<=signed(MULTS_5_1(5)(PRECISION-1 downto 0))+signed(MULTS_5_2(5)(PRECISION-1 downto 0));
			MULTS_6_1(6)<=signed(MULTS_5_1(6)(PRECISION-1 downto 0))+signed(MULTS_5_2(6)(PRECISION-1 downto 0));
			MULTS_6_1(7)<=signed(MULTS_5_1(7)(PRECISION-1 downto 0))+signed(MULTS_5_2(7)(PRECISION-1 downto 0));
			MULTS_6_1(8)<=signed(MULTS_5_1(8)(PRECISION-1 downto 0))+signed(MULTS_5_2(8)(PRECISION-1 downto 0));
			MULTS_6_1(9)<=signed(MULTS_5_1(9)(PRECISION-1 downto 0))+signed(MULTS_5_2(9)(PRECISION-1 downto 0));



                         EN_SUM_MULT_7<='1';
		end if;


		------------------------- Enable NEXT STATGE MULTS START -----------------------

		if EN_SUM_MULT_7 = '1' then
			------------------------------------STAGE-7--------------------------------------
			MULTS_7_1(0)<=signed(MULTS_6_1(0)(PRECISION-1 downto 0))+signed(MULTS_6_2(0)(PRECISION-1 downto 0));
			MULTS_7_1(1)<=signed(MULTS_6_1(1)(PRECISION-1 downto 0))+signed(MULTS_6_2(1)(PRECISION-1 downto 0));
			MULTS_7_1(2)<=signed(MULTS_6_1(2)(PRECISION-1 downto 0))+signed(MULTS_6_2(2)(PRECISION-1 downto 0));
			MULTS_7_1(3)<=signed(MULTS_6_1(3)(PRECISION-1 downto 0))+signed(MULTS_6_2(3)(PRECISION-1 downto 0));
			MULTS_7_1(4)<=signed(MULTS_6_1(4)(PRECISION-1 downto 0))+signed(MULTS_6_2(4)(PRECISION-1 downto 0));
			MULTS_7_1(5)<=signed(MULTS_6_1(5)(PRECISION-1 downto 0))+signed(MULTS_6_2(5)(PRECISION-1 downto 0));
			MULTS_7_1(6)<=signed(MULTS_6_1(6)(PRECISION-1 downto 0))+signed(MULTS_6_2(6)(PRECISION-1 downto 0));
			MULTS_7_1(7)<=signed(MULTS_6_1(7)(PRECISION-1 downto 0))+signed(MULTS_6_2(7)(PRECISION-1 downto 0));
			MULTS_7_1(8)<=signed(MULTS_6_1(8)(PRECISION-1 downto 0))+signed(MULTS_6_2(8)(PRECISION-1 downto 0));
			MULTS_7_1(9)<=signed(MULTS_6_1(9)(PRECISION-1 downto 0))+signed(MULTS_6_2(9)(PRECISION-1 downto 0));



                        Enable_BIAS<='1';
		end if;


		------------------------------------STAGE-BIAS--------------------------------------
		if Enable_BIAS = '1' then

			BIAS_1<=(signed(BIAS_VAL_1)+ signed(MULTS_7_1(0)(PRECISION-1 downto 0)));
			BIAS_2<=(signed(BIAS_VAL_2)+ signed(MULTS_7_1(1)(PRECISION-1 downto 0)));
			BIAS_3<=(signed(BIAS_VAL_3)+ signed(MULTS_7_1(2)(PRECISION-1 downto 0)));
			BIAS_4<=(signed(BIAS_VAL_4)+ signed(MULTS_7_1(3)(PRECISION-1 downto 0)));
			BIAS_5<=(signed(BIAS_VAL_5)+ signed(MULTS_7_1(4)(PRECISION-1 downto 0)));
			BIAS_6<=(signed(BIAS_VAL_6)+ signed(MULTS_7_1(5)(PRECISION-1 downto 0)));
			BIAS_7<=(signed(BIAS_VAL_7)+ signed(MULTS_7_1(6)(PRECISION-1 downto 0)));
			BIAS_8<=(signed(BIAS_VAL_8)+ signed(MULTS_7_1(7)(PRECISION-1 downto 0)));
			BIAS_9<=(signed(BIAS_VAL_9)+ signed(MULTS_7_1(8)(PRECISION-1 downto 0)));
			BIAS_10<=(signed(BIAS_VAL_10)+ signed(MULTS_7_1(9)(PRECISION-1 downto 0)));

			Enable_ReLU<='1';
			
		end if;

		if SIG_STRIDE>1 and Enable_ReLU='1' then
                 SIG_STRIDE<=SIG_STRIDE-1; end if;

	if  Enable_ReLU='1' then
		if VALID_NXTLYR_PIX<VALID_LOCAL_PIX and SIG_STRIDE>(STRIDE-1) then

			if BIAS_1>0 then
			ReLU_1<=BIAS_1;
			DOUT_BUF_1_7<=std_logic_vector(BIAS_1);
			else
			ReLU_1<= (others => '0');
			DOUT_BUF_1_7<=(others => '0');
			end if;
			if BIAS_2>0 then
			ReLU_2<=BIAS_2;
			DOUT_BUF_2_7<=std_logic_vector(BIAS_2);
			else
			ReLU_2<= (others => '0');
			DOUT_BUF_2_7<=(others => '0');
			end if;
			if BIAS_3>0 then
			ReLU_3<=BIAS_3;
			DOUT_BUF_3_7<=std_logic_vector(BIAS_3);
			else
			ReLU_3<= (others => '0');
			DOUT_BUF_3_7<=(others => '0');
			end if;
			if BIAS_4>0 then
			ReLU_4<=BIAS_4;
			DOUT_BUF_4_7<=std_logic_vector(BIAS_4);
			else
			ReLU_4<= (others => '0');
			DOUT_BUF_4_7<=(others => '0');
			end if;
			if BIAS_5>0 then
			ReLU_5<=BIAS_5;
			DOUT_BUF_5_7<=std_logic_vector(BIAS_5);
			else
			ReLU_5<= (others => '0');
			DOUT_BUF_5_7<=(others => '0');
			end if;
			if BIAS_6>0 then
			ReLU_6<=BIAS_6;
			DOUT_BUF_6_7<=std_logic_vector(BIAS_6);
			else
			ReLU_6<= (others => '0');
			DOUT_BUF_6_7<=(others => '0');
			end if;
			if BIAS_7>0 then
			ReLU_7<=BIAS_7;
			DOUT_BUF_7_7<=std_logic_vector(BIAS_7);
			else
			ReLU_7<= (others => '0');
			DOUT_BUF_7_7<=(others => '0');
			end if;
			if BIAS_8>0 then
			ReLU_8<=BIAS_8;
			DOUT_BUF_8_7<=std_logic_vector(BIAS_8);
			else
			ReLU_8<= (others => '0');
			DOUT_BUF_8_7<=(others => '0');
			end if;
			if BIAS_9>0 then
			ReLU_9<=BIAS_9;
			DOUT_BUF_9_7<=std_logic_vector(BIAS_9);
			else
			ReLU_9<= (others => '0');
			DOUT_BUF_9_7<=(others => '0');
			end if;
			if BIAS_10>0 then
			ReLU_10<=BIAS_10;
			DOUT_BUF_10_7<=std_logic_vector(BIAS_10);
			else
			ReLU_10<= (others => '0');
			DOUT_BUF_10_7<=(others => '0');
			end if;

			EN_NXT_LYR_7<='1';FRST_TIM_EN_7<='1';
			OUT_PIXEL_COUNT<=OUT_PIXEL_COUNT+1;
		else
                       EN_NXT_LYR_7<='0';
                       DOUT_BUF_1_7<=(others => '0');
                       DOUT_BUF_2_7<=(others => '0');
                       DOUT_BUF_3_7<=(others => '0');
                       DOUT_BUF_4_7<=(others => '0');
                       DOUT_BUF_5_7<=(others => '0');
                       DOUT_BUF_6_7<=(others => '0');
                       DOUT_BUF_7_7<=(others => '0');
                       DOUT_BUF_8_7<=(others => '0');
                       DOUT_BUF_9_7<=(others => '0');
                       DOUT_BUF_10_7<=(others => '0');

		end if; -- VALIDPIXELS

		if VALID_NXTLYR_PIX=((VALID_LOCAL_PIX*STRIDE)-1) then VALID_NXTLYR_PIX<=0;SIG_STRIDE<=STRIDE;   -- reset sride and valid pixels
		else VALID_NXTLYR_PIX<=VALID_NXTLYR_PIX+1;end if; 

	end if;  --ReLU
elsif OUT_PIXEL_COUNT>=VALID_CYCLES  then INTERNAL_RST<='1';SIG_STRIDE<=STRIDE;EN_NXT_LYR_7<='1';  -- order is very important
else  EN_NXT_LYR_7<='0';-- In case stream stopped

end if; -- end enable 
end if; -- for RST	
end if; -- rising edge
end process LAYER_7;

DOUT_1_7<=DOUT_BUF_1_7;
DOUT_2_7<=DOUT_BUF_2_7;
DOUT_3_7<=DOUT_BUF_3_7;
DOUT_4_7<=DOUT_BUF_4_7;
DOUT_5_7<=DOUT_BUF_5_7;
DOUT_6_7<=DOUT_BUF_6_7;
DOUT_7_7<=DOUT_BUF_7_7;
DOUT_8_7<=DOUT_BUF_8_7;
DOUT_9_7<=DOUT_BUF_9_7;
DOUT_10_7<=DOUT_BUF_10_7;

end Behavioral;
------------------------------ ARCHITECTURE DECLARATION - END---------------------------------------------

